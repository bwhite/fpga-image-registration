/home/brandyn/fpga-image-registration/modules/./smooth_stage/smooth_address_selector.vhd