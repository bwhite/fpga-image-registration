/home/brandyn/fpga-image-registration/modules/./make_h_matrix/make_h_matrix.vhd