/home/brandyn/fpga-image-registration/modules/./make_affine_homography/make_affine_homography.vhd