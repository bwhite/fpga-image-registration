/home/brandyn/fpga-image-registration/modules/./registration_stage/registration_stage.vhd