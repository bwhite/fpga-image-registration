LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
ENTITY gauss_elimT0_tb IS
PORT(
  CLK : IN STD_LOGIC;
  RST : IN STD_LOGIC;
  DONE : OUT STD_LOGIC;
  FAIL : OUT STD_LOGIC;
  FAIL_NUM : OUT STD_LOGIC_VECTOR(10 DOWNTO 0));
END gauss_elimT0_tb;
ARCHITECTURE behavior OF gauss_elimT0_tb IS
  COMPONENT gauss_elim
  PORT(
    CLK : IN STD_LOGIC;
    RST : IN STD_LOGIC;
    INPUT_LOAD : IN STD_LOGIC;
    A_0_0 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_0_1 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_0_2 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_0_3 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_0_4 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_0_5 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_1_0 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_1_1 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_1_2 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_1_3 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_1_4 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_1_5 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_2_0 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_2_1 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_2_2 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_2_3 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_2_4 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_2_5 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_3_0 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_3_1 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_3_2 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_3_3 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_3_4 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_3_5 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_4_0 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_4_1 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_4_2 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_4_3 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_4_4 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_4_5 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_5_0 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_5_1 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_5_2 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_5_3 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_5_4 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_5_5 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    B_0 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    B_1 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    B_2 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    B_3 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    B_4 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    B_5 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    X_0 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    X_1 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    X_2 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    X_3 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    X_4 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    X_5 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    OUTPUT_VALID : OUT STD_LOGIC);
  END COMPONENT;
  SIGNAL uut_rst_wire, uut_rst : STD_LOGIC;
  SIGNAL state : STD_LOGIC_VECTOR(10 DOWNTO 0);
  -- UUT Input
  SIGNAL uut_input_load : STD_LOGIC;
  SIGNAL uut_a_0_0, uut_a_0_1, uut_a_0_2, uut_a_0_3, uut_a_0_4, uut_a_0_5, uut_a_1_0, uut_a_1_1, uut_a_1_2, uut_a_1_3, uut_a_1_4, uut_a_1_5, uut_a_2_0, uut_a_2_1, uut_a_2_2, uut_a_2_3, uut_a_2_4, uut_a_2_5, uut_a_3_0, uut_a_3_1, uut_a_3_2, uut_a_3_3, uut_a_3_4, uut_a_3_5, uut_a_4_0, uut_a_4_1, uut_a_4_2, uut_a_4_3, uut_a_4_4, uut_a_4_5, uut_a_5_0, uut_a_5_1, uut_a_5_2, uut_a_5_3, uut_a_5_4, uut_a_5_5, uut_b_0, uut_b_1, uut_b_2, uut_b_3, uut_b_4, uut_b_5 : STD_LOGIC_VECTOR(26 DOWNTO 0);
  -- UUT Output
  SIGNAL uut_output_valid : STD_LOGIC;
  SIGNAL uut_x_0, uut_x_1, uut_x_2, uut_x_3, uut_x_4, uut_x_5 : STD_LOGIC_VECTOR(26 DOWNTO 0);
BEGIN
  uut_rst_wire <= RST OR uut_rst;
  uut :  gauss_elim PORT MAP (
    CLK => CLK,
    RST => uut_rst_wire,
    INPUT_LOAD => uut_input_load,
    A_0_0 => uut_a_0_0,
    A_0_1 => uut_a_0_1,
    A_0_2 => uut_a_0_2,
    A_0_3 => uut_a_0_3,
    A_0_4 => uut_a_0_4,
    A_0_5 => uut_a_0_5,
    A_1_0 => uut_a_1_0,
    A_1_1 => uut_a_1_1,
    A_1_2 => uut_a_1_2,
    A_1_3 => uut_a_1_3,
    A_1_4 => uut_a_1_4,
    A_1_5 => uut_a_1_5,
    A_2_0 => uut_a_2_0,
    A_2_1 => uut_a_2_1,
    A_2_2 => uut_a_2_2,
    A_2_3 => uut_a_2_3,
    A_2_4 => uut_a_2_4,
    A_2_5 => uut_a_2_5,
    A_3_0 => uut_a_3_0,
    A_3_1 => uut_a_3_1,
    A_3_2 => uut_a_3_2,
    A_3_3 => uut_a_3_3,
    A_3_4 => uut_a_3_4,
    A_3_5 => uut_a_3_5,
    A_4_0 => uut_a_4_0,
    A_4_1 => uut_a_4_1,
    A_4_2 => uut_a_4_2,
    A_4_3 => uut_a_4_3,
    A_4_4 => uut_a_4_4,
    A_4_5 => uut_a_4_5,
    A_5_0 => uut_a_5_0,
    A_5_1 => uut_a_5_1,
    A_5_2 => uut_a_5_2,
    A_5_3 => uut_a_5_3,
    A_5_4 => uut_a_5_4,
    A_5_5 => uut_a_5_5,
    B_0 => uut_b_0,
    B_1 => uut_b_1,
    B_2 => uut_b_2,
    B_3 => uut_b_3,
    B_4 => uut_b_4,
    B_5 => uut_b_5,
    X_0 => uut_x_0,
    X_1 => uut_x_1,
    X_2 => uut_x_2,
    X_3 => uut_x_3,
    X_4 => uut_x_4,
    X_5 => uut_x_5,
    OUTPUT_VALID => uut_output_valid
  );
  PROCESS (CLK) IS
  BEGIN
    IF CLK'event AND CLK='1' THEN
      IF RST='1' THEN
        DONE <= '0';
        FAIL <= '0';
        uut_rst <= '1';
        FAIL_NUM <= (OTHERS => '0');
        state <= (OTHERS => '0');
      ELSE
        CASE state IS
          WHEN "00000000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000000001";
            uut_rst <= '0';
          WHEN "00000000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000000010";
            uut_rst <= '0';
          WHEN "00000000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000000011";
            uut_rst <= '0';
          WHEN "00000000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000000100";
            uut_rst <= '0';
          WHEN "00000000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000000101";
            uut_rst <= '0';
          WHEN "00000000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000000110";
            uut_rst <= '0';
          WHEN "00000000110" =>
            uut_input_load <= '1';
            uut_a_0_0 <= "000000000011000011010110100";
            uut_a_0_1 <= "000000001100111111000011100";
            uut_a_0_2 <= "000000111001100101001111000";
            uut_a_0_3 <= "000000000000000010001010010";
            uut_a_0_4 <= "000000000111100110101010100";
            uut_a_0_5 <= "111111111101000110011001000";
            uut_a_1_0 <= "000000000000000110011111100";
            uut_a_1_1 <= "000000100010110101001001111";
            uut_a_1_2 <= "000000000110100011000110110";
            uut_a_1_3 <= "000000000000000011110011010";
            uut_a_1_4 <= "111111111111110101011011101";
            uut_a_1_5 <= "000000000000010010011110001";
            uut_a_2_0 <= "000000000000011100110010100";
            uut_a_2_1 <= "000000000110100011000110110";
            uut_a_2_2 <= "000000010011101111110011100";
            uut_a_2_3 <= "111111111111111110100011001";
            uut_a_2_4 <= "000000000000010010011110001";
            uut_a_2_5 <= "111111111110101101111000110";
            uut_a_3_0 <= "000000000000000010001010010";
            uut_a_3_1 <= "000000000111100110101010100";
            uut_a_3_2 <= "111111111101000110011001000";
            uut_a_3_3 <= "000000000100001110101100001";
            uut_a_3_4 <= "000001101101010011010000101";
            uut_a_3_5 <= "000000011110111111111010000";
            uut_a_4_0 <= "000000000000000011110011010";
            uut_a_4_1 <= "111111111111110101011011101";
            uut_a_4_2 <= "000000000000010010011110001";
            uut_a_4_3 <= "000000000000110110101001101";
            uut_a_4_4 <= "000001000000011100000111000";
            uut_a_4_5 <= "000000000011100110111011111";
            uut_a_5_0 <= "111111111111111110100011001";
            uut_a_5_1 <= "000000000000010010011110001";
            uut_a_5_2 <= "111111111110101101111000110";
            uut_a_5_3 <= "000000000000001111011111111";
            uut_a_5_4 <= "000000000011100110111011111";
            uut_a_5_5 <= "000000010101101100011000110";
            state <= "00000000111";
            uut_rst <= '0';
          WHEN "00000000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000001000";
            uut_rst <= '0';
          WHEN "00000001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000001001";
            uut_rst <= '0';
          WHEN "00000001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000001010";
            uut_rst <= '0';
          WHEN "00000001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000001011";
            uut_rst <= '0';
          WHEN "00000001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000001100";
            uut_rst <= '0';
          WHEN "00000001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000001101";
            uut_rst <= '0';
          WHEN "00000001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000001110";
            uut_rst <= '0';
          WHEN "00000001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000001111";
            uut_rst <= '0';
          WHEN "00000001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000010000";
            uut_rst <= '0';
          WHEN "00000010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000010001";
            uut_rst <= '0';
          WHEN "00000010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000010010";
            uut_rst <= '0';
          WHEN "00000010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000010011";
            uut_rst <= '0';
          WHEN "00000010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000010100";
            uut_rst <= '0';
          WHEN "00000010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000010101";
            uut_rst <= '0';
          WHEN "00000010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000010110";
            uut_rst <= '0';
          WHEN "00000010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000010111";
            uut_rst <= '0';
          WHEN "00000010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000011000";
            uut_rst <= '0';
          WHEN "00000011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000011001";
            uut_rst <= '0';
          WHEN "00000011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000011010";
            uut_rst <= '0';
          WHEN "00000011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000011011";
            uut_rst <= '0';
          WHEN "00000011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000011100";
            uut_rst <= '0';
          WHEN "00000011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000011101";
            uut_rst <= '0';
          WHEN "00000011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000011110";
            uut_rst <= '0';
          WHEN "00000011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000011111";
            uut_rst <= '0';
          WHEN "00000011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000100000";
            uut_rst <= '0';
          WHEN "00000100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000100001";
            uut_rst <= '0';
          WHEN "00000100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000100010";
            uut_rst <= '0';
          WHEN "00000100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000100011";
            uut_rst <= '0';
          WHEN "00000100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000100100";
            uut_rst <= '0';
          WHEN "00000100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000100101";
            uut_rst <= '0';
          WHEN "00000100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000100110";
            uut_rst <= '0';
          WHEN "00000100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000100111";
            uut_rst <= '0';
          WHEN "00000100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000101000";
            uut_rst <= '0';
          WHEN "00000101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000101001";
            uut_rst <= '0';
          WHEN "00000101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000101010";
            uut_rst <= '0';
          WHEN "00000101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000101011";
            uut_rst <= '0';
          WHEN "00000101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000101100";
            uut_rst <= '0';
          WHEN "00000101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000101101";
            uut_rst <= '0';
          WHEN "00000101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000101110";
            uut_rst <= '0';
          WHEN "00000101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000101111";
            uut_rst <= '0';
          WHEN "00000101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000110000";
            uut_rst <= '0';
          WHEN "00000110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000110001";
            uut_rst <= '0';
          WHEN "00000110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000110010";
            uut_rst <= '0';
          WHEN "00000110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000110011";
            uut_rst <= '0';
          WHEN "00000110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000110100";
            uut_rst <= '0';
          WHEN "00000110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000110101";
            uut_rst <= '0';
          WHEN "00000110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000110110";
            uut_rst <= '0';
          WHEN "00000110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000110111";
            uut_rst <= '0';
          WHEN "00000110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000111000";
            uut_rst <= '0';
          WHEN "00000111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000111001";
            uut_rst <= '0';
          WHEN "00000111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000111010";
            uut_rst <= '0';
          WHEN "00000111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000111011";
            uut_rst <= '0';
          WHEN "00000111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000111100";
            uut_rst <= '0';
          WHEN "00000111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000111101";
            uut_rst <= '0';
          WHEN "00000111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000111110";
            uut_rst <= '0';
          WHEN "00000111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00000111111";
            uut_rst <= '0';
          WHEN "00000111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001000000";
            uut_rst <= '0';
          WHEN "00001000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001000001";
            uut_rst <= '0';
          WHEN "00001000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001000010";
            uut_rst <= '0';
          WHEN "00001000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001000011";
            uut_rst <= '0';
          WHEN "00001000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001000100";
            uut_rst <= '0';
          WHEN "00001000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001000101";
            uut_rst <= '0';
          WHEN "00001000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001000110";
            uut_rst <= '0';
          WHEN "00001000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001000111";
            uut_rst <= '0';
          WHEN "00001000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001001000";
            uut_rst <= '0';
          WHEN "00001001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001001001";
            uut_rst <= '0';
          WHEN "00001001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001001010";
            uut_rst <= '0';
          WHEN "00001001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001001011";
            uut_rst <= '0';
          WHEN "00001001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001001100";
            uut_rst <= '0';
          WHEN "00001001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001001101";
            uut_rst <= '0';
          WHEN "00001001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001001110";
            uut_rst <= '0';
          WHEN "00001001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001001111";
            uut_rst <= '0';
          WHEN "00001001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001010000";
            uut_rst <= '0';
          WHEN "00001010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001010001";
            uut_rst <= '0';
          WHEN "00001010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001010010";
            uut_rst <= '0';
          WHEN "00001010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001010011";
            uut_rst <= '0';
          WHEN "00001010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001010100";
            uut_rst <= '0';
          WHEN "00001010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001010101";
            uut_rst <= '0';
          WHEN "00001010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001010110";
            uut_rst <= '0';
          WHEN "00001010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001010111";
            uut_rst <= '0';
          WHEN "00001010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001011000";
            uut_rst <= '0';
          WHEN "00001011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001011001";
            uut_rst <= '0';
          WHEN "00001011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001011010";
            uut_rst <= '0';
          WHEN "00001011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001011011";
            uut_rst <= '0';
          WHEN "00001011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001011100";
            uut_rst <= '0';
          WHEN "00001011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001011101";
            uut_rst <= '0';
          WHEN "00001011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001011110";
            uut_rst <= '0';
          WHEN "00001011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001011111";
            uut_rst <= '0';
          WHEN "00001011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001100000";
            uut_rst <= '0';
          WHEN "00001100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001100001";
            uut_rst <= '0';
          WHEN "00001100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001100010";
            uut_rst <= '0';
          WHEN "00001100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001100011";
            uut_rst <= '0';
          WHEN "00001100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001100100";
            uut_rst <= '0';
          WHEN "00001100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001100101";
            uut_rst <= '0';
          WHEN "00001100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001100110";
            uut_rst <= '0';
          WHEN "00001100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001100111";
            uut_rst <= '0';
          WHEN "00001100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001101000";
            uut_rst <= '0';
          WHEN "00001101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001101001";
            uut_rst <= '0';
          WHEN "00001101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001101010";
            uut_rst <= '0';
          WHEN "00001101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001101011";
            uut_rst <= '0';
          WHEN "00001101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001101100";
            uut_rst <= '0';
          WHEN "00001101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001101101";
            uut_rst <= '0';
          WHEN "00001101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001101110";
            uut_rst <= '0';
          WHEN "00001101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001101111";
            uut_rst <= '0';
          WHEN "00001101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001110000";
            uut_rst <= '0';
          WHEN "00001110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001110001";
            uut_rst <= '0';
          WHEN "00001110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001110010";
            uut_rst <= '0';
          WHEN "00001110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001110011";
            uut_rst <= '0';
          WHEN "00001110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001110100";
            uut_rst <= '0';
          WHEN "00001110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001110101";
            uut_rst <= '0';
          WHEN "00001110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001110110";
            uut_rst <= '0';
          WHEN "00001110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001110111";
            uut_rst <= '0';
          WHEN "00001110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001111000";
            uut_rst <= '0';
          WHEN "00001111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001111001";
            uut_rst <= '0';
          WHEN "00001111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001111010";
            uut_rst <= '0';
          WHEN "00001111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001111011";
            uut_rst <= '0';
          WHEN "00001111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001111100";
            uut_rst <= '0';
          WHEN "00001111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001111101";
            uut_rst <= '0';
          WHEN "00001111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001111110";
            uut_rst <= '0';
          WHEN "00001111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00001111111";
            uut_rst <= '0';
          WHEN "00001111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010000000";
            uut_rst <= '0';
          WHEN "00010000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010000001";
            uut_rst <= '0';
          WHEN "00010000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010000010";
            uut_rst <= '0';
          WHEN "00010000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010000011";
            uut_rst <= '0';
          WHEN "00010000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010000100";
            uut_rst <= '0';
          WHEN "00010000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010000101";
            uut_rst <= '0';
          WHEN "00010000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010000110";
            uut_rst <= '0';
          WHEN "00010000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010000111";
            uut_rst <= '0';
          WHEN "00010000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010001000";
            uut_rst <= '0';
          WHEN "00010001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010001001";
            uut_rst <= '0';
          WHEN "00010001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010001010";
            uut_rst <= '0';
          WHEN "00010001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010001011";
            uut_rst <= '0';
          WHEN "00010001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010001100";
            uut_rst <= '0';
          WHEN "00010001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010001101";
            uut_rst <= '0';
          WHEN "00010001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010001110";
            uut_rst <= '0';
          WHEN "00010001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010001111";
            uut_rst <= '0';
          WHEN "00010001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010010000";
            uut_rst <= '0';
          WHEN "00010010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010010001";
            uut_rst <= '0';
          WHEN "00010010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010010010";
            uut_rst <= '0';
          WHEN "00010010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010010011";
            uut_rst <= '0';
          WHEN "00010010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010010100";
            uut_rst <= '0';
          WHEN "00010010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010010101";
            uut_rst <= '0';
          WHEN "00010010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010010110";
            uut_rst <= '0';
          WHEN "00010010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010010111";
            uut_rst <= '0';
          WHEN "00010010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010011000";
            uut_rst <= '0';
          WHEN "00010011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010011001";
            uut_rst <= '0';
          WHEN "00010011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010011010";
            uut_rst <= '0';
          WHEN "00010011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010011011";
            uut_rst <= '0';
          WHEN "00010011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010011100";
            uut_rst <= '0';
          WHEN "00010011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010011101";
            uut_rst <= '0';
          WHEN "00010011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010011110";
            uut_rst <= '0';
          WHEN "00010011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010011111";
            uut_rst <= '0';
          WHEN "00010011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010100000";
            uut_rst <= '0';
          WHEN "00010100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010100001";
            uut_rst <= '0';
          WHEN "00010100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010100010";
            uut_rst <= '0';
          WHEN "00010100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010100011";
            uut_rst <= '0';
          WHEN "00010100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010100100";
            uut_rst <= '0';
          WHEN "00010100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010100101";
            uut_rst <= '0';
          WHEN "00010100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010100110";
            uut_rst <= '0';
          WHEN "00010100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010100111";
            uut_rst <= '0';
          WHEN "00010100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010101000";
            uut_rst <= '0';
          WHEN "00010101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010101001";
            uut_rst <= '0';
          WHEN "00010101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010101010";
            uut_rst <= '0';
          WHEN "00010101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010101011";
            uut_rst <= '0';
          WHEN "00010101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010101100";
            uut_rst <= '0';
          WHEN "00010101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010101101";
            uut_rst <= '0';
          WHEN "00010101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010101110";
            uut_rst <= '0';
          WHEN "00010101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010101111";
            uut_rst <= '0';
          WHEN "00010101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010110000";
            uut_rst <= '0';
          WHEN "00010110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010110001";
            uut_rst <= '0';
          WHEN "00010110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010110010";
            uut_rst <= '0';
          WHEN "00010110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010110011";
            uut_rst <= '0';
          WHEN "00010110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010110100";
            uut_rst <= '0';
          WHEN "00010110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010110101";
            uut_rst <= '0';
          WHEN "00010110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010110110";
            uut_rst <= '0';
          WHEN "00010110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010110111";
            uut_rst <= '0';
          WHEN "00010110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010111000";
            uut_rst <= '0';
          WHEN "00010111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010111001";
            uut_rst <= '0';
          WHEN "00010111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010111010";
            uut_rst <= '0';
          WHEN "00010111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010111011";
            uut_rst <= '0';
          WHEN "00010111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010111100";
            uut_rst <= '0';
          WHEN "00010111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010111101";
            uut_rst <= '0';
          WHEN "00010111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010111110";
            uut_rst <= '0';
          WHEN "00010111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00010111111";
            uut_rst <= '0';
          WHEN "00010111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011000000";
            uut_rst <= '0';
          WHEN "00011000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011000001";
            uut_rst <= '0';
          WHEN "00011000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011000010";
            uut_rst <= '0';
          WHEN "00011000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011000011";
            uut_rst <= '0';
          WHEN "00011000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011000100";
            uut_rst <= '0';
          WHEN "00011000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011000101";
            uut_rst <= '0';
          WHEN "00011000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011000110";
            uut_rst <= '0';
          WHEN "00011000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011000111";
            uut_rst <= '0';
          WHEN "00011000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011001000";
            uut_rst <= '0';
          WHEN "00011001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011001001";
            uut_rst <= '0';
          WHEN "00011001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011001010";
            uut_rst <= '0';
          WHEN "00011001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011001011";
            uut_rst <= '0';
          WHEN "00011001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011001100";
            uut_rst <= '0';
          WHEN "00011001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011001101";
            uut_rst <= '0';
          WHEN "00011001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011001110";
            uut_rst <= '0';
          WHEN "00011001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011001111";
            uut_rst <= '0';
          WHEN "00011001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011010000";
            uut_rst <= '0';
          WHEN "00011010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011010001";
            uut_rst <= '0';
          WHEN "00011010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011010010";
            uut_rst <= '0';
          WHEN "00011010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011010011";
            uut_rst <= '0';
          WHEN "00011010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011010100";
            uut_rst <= '0';
          WHEN "00011010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011010101";
            uut_rst <= '0';
          WHEN "00011010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011010110";
            uut_rst <= '0';
          WHEN "00011010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011010111";
            uut_rst <= '0';
          WHEN "00011010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011011000";
            uut_rst <= '0';
          WHEN "00011011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011011001";
            uut_rst <= '0';
          WHEN "00011011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011011010";
            uut_rst <= '0';
          WHEN "00011011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011011011";
            uut_rst <= '0';
          WHEN "00011011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011011100";
            uut_rst <= '0';
          WHEN "00011011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011011101";
            uut_rst <= '0';
          WHEN "00011011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011011110";
            uut_rst <= '0';
          WHEN "00011011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011011111";
            uut_rst <= '0';
          WHEN "00011011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011100000";
            uut_rst <= '0';
          WHEN "00011100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011100001";
            uut_rst <= '0';
          WHEN "00011100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011100010";
            uut_rst <= '0';
          WHEN "00011100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011100011";
            uut_rst <= '0';
          WHEN "00011100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011100100";
            uut_rst <= '0';
          WHEN "00011100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011100101";
            uut_rst <= '0';
          WHEN "00011100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011100110";
            uut_rst <= '0';
          WHEN "00011100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011100111";
            uut_rst <= '0';
          WHEN "00011100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011101000";
            uut_rst <= '0';
          WHEN "00011101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011101001";
            uut_rst <= '0';
          WHEN "00011101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011101010";
            uut_rst <= '0';
          WHEN "00011101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011101011";
            uut_rst <= '0';
          WHEN "00011101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011101100";
            uut_rst <= '0';
          WHEN "00011101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011101101";
            uut_rst <= '0';
          WHEN "00011101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011101110";
            uut_rst <= '0';
          WHEN "00011101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011101111";
            uut_rst <= '0';
          WHEN "00011101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011110000";
            uut_rst <= '0';
          WHEN "00011110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011110001";
            uut_rst <= '0';
          WHEN "00011110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011110010";
            uut_rst <= '0';
          WHEN "00011110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011110011";
            uut_rst <= '0';
          WHEN "00011110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011110100";
            uut_rst <= '0';
          WHEN "00011110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011110101";
            uut_rst <= '0';
          WHEN "00011110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011110110";
            uut_rst <= '0';
          WHEN "00011110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011110111";
            uut_rst <= '0';
          WHEN "00011110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011111000";
            uut_rst <= '0';
          WHEN "00011111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011111001";
            uut_rst <= '0';
          WHEN "00011111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011111010";
            uut_rst <= '0';
          WHEN "00011111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011111011";
            uut_rst <= '0';
          WHEN "00011111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011111100";
            uut_rst <= '0';
          WHEN "00011111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011111101";
            uut_rst <= '0';
          WHEN "00011111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011111110";
            uut_rst <= '0';
          WHEN "00011111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00011111111";
            uut_rst <= '0';
          WHEN "00011111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100000000";
            uut_rst <= '0';
          WHEN "00100000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100000001";
            uut_rst <= '0';
          WHEN "00100000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100000010";
            uut_rst <= '0';
          WHEN "00100000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100000011";
            uut_rst <= '0';
          WHEN "00100000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100000100";
            uut_rst <= '0';
          WHEN "00100000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100000101";
            uut_rst <= '0';
          WHEN "00100000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100000110";
            uut_rst <= '0';
          WHEN "00100000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100000111";
            uut_rst <= '0';
          WHEN "00100000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100001000";
            uut_rst <= '0';
          WHEN "00100001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100001001";
            uut_rst <= '0';
          WHEN "00100001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100001010";
            uut_rst <= '0';
          WHEN "00100001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100001011";
            uut_rst <= '0';
          WHEN "00100001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100001100";
            uut_rst <= '0';
          WHEN "00100001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100001101";
            uut_rst <= '0';
          WHEN "00100001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100001110";
            uut_rst <= '0';
          WHEN "00100001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100001111";
            uut_rst <= '0';
          WHEN "00100001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100010000";
            uut_rst <= '0';
          WHEN "00100010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100010001";
            uut_rst <= '0';
          WHEN "00100010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100010010";
            uut_rst <= '0';
          WHEN "00100010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100010011";
            uut_rst <= '0';
          WHEN "00100010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100010100";
            uut_rst <= '0';
          WHEN "00100010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100010101";
            uut_rst <= '0';
          WHEN "00100010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100010110";
            uut_rst <= '0';
          WHEN "00100010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100010111";
            uut_rst <= '0';
          WHEN "00100010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100011000";
            uut_rst <= '0';
          WHEN "00100011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100011001";
            uut_rst <= '0';
          WHEN "00100011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100011010";
            uut_rst <= '0';
          WHEN "00100011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100011011";
            uut_rst <= '0';
          WHEN "00100011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100011100";
            uut_rst <= '0';
          WHEN "00100011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100011101";
            uut_rst <= '0';
          WHEN "00100011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100011110";
            uut_rst <= '0';
          WHEN "00100011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100011111";
            uut_rst <= '0';
          WHEN "00100011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100100000";
            uut_rst <= '0';
          WHEN "00100100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100100001";
            uut_rst <= '0';
          WHEN "00100100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100100010";
            uut_rst <= '0';
          WHEN "00100100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100100011";
            uut_rst <= '0';
          WHEN "00100100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100100100";
            uut_rst <= '0';
          WHEN "00100100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100100101";
            uut_rst <= '0';
          WHEN "00100100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100100110";
            uut_rst <= '0';
          WHEN "00100100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100100111";
            uut_rst <= '0';
          WHEN "00100100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100101000";
            uut_rst <= '0';
          WHEN "00100101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100101001";
            uut_rst <= '0';
          WHEN "00100101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100101010";
            uut_rst <= '0';
          WHEN "00100101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100101011";
            uut_rst <= '0';
          WHEN "00100101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100101100";
            uut_rst <= '0';
          WHEN "00100101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100101101";
            uut_rst <= '0';
          WHEN "00100101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100101110";
            uut_rst <= '0';
          WHEN "00100101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100101111";
            uut_rst <= '0';
          WHEN "00100101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100110000";
            uut_rst <= '0';
          WHEN "00100110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100110001";
            uut_rst <= '0';
          WHEN "00100110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100110010";
            uut_rst <= '0';
          WHEN "00100110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100110011";
            uut_rst <= '0';
          WHEN "00100110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100110100";
            uut_rst <= '0';
          WHEN "00100110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100110101";
            uut_rst <= '0';
          WHEN "00100110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100110110";
            uut_rst <= '0';
          WHEN "00100110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100110111";
            uut_rst <= '0';
          WHEN "00100110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100111000";
            uut_rst <= '0';
          WHEN "00100111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100111001";
            uut_rst <= '0';
          WHEN "00100111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100111010";
            uut_rst <= '0';
          WHEN "00100111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100111011";
            uut_rst <= '0';
          WHEN "00100111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100111100";
            uut_rst <= '0';
          WHEN "00100111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100111101";
            uut_rst <= '0';
          WHEN "00100111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100111110";
            uut_rst <= '0';
          WHEN "00100111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00100111111";
            uut_rst <= '0';
          WHEN "00100111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101000000";
            uut_rst <= '0';
          WHEN "00101000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101000001";
            uut_rst <= '0';
          WHEN "00101000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101000010";
            uut_rst <= '0';
          WHEN "00101000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101000011";
            uut_rst <= '0';
          WHEN "00101000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101000100";
            uut_rst <= '0';
          WHEN "00101000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101000101";
            uut_rst <= '0';
          WHEN "00101000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101000110";
            uut_rst <= '0';
          WHEN "00101000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101000111";
            uut_rst <= '0';
          WHEN "00101000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101001000";
            uut_rst <= '0';
          WHEN "00101001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101001001";
            uut_rst <= '0';
          WHEN "00101001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101001010";
            uut_rst <= '0';
          WHEN "00101001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101001011";
            uut_rst <= '0';
          WHEN "00101001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101001100";
            uut_rst <= '0';
          WHEN "00101001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101001101";
            uut_rst <= '0';
          WHEN "00101001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101001110";
            uut_rst <= '0';
          WHEN "00101001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101001111";
            uut_rst <= '0';
          WHEN "00101001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101010000";
            uut_rst <= '0';
          WHEN "00101010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101010001";
            uut_rst <= '0';
          WHEN "00101010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101010010";
            uut_rst <= '0';
          WHEN "00101010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101010011";
            uut_rst <= '0';
          WHEN "00101010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101010100";
            uut_rst <= '0';
          WHEN "00101010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101010101";
            uut_rst <= '0';
          WHEN "00101010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101010110";
            uut_rst <= '0';
          WHEN "00101010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101010111";
            uut_rst <= '0';
          WHEN "00101010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101011000";
            uut_rst <= '0';
          WHEN "00101011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101011001";
            uut_rst <= '0';
          WHEN "00101011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101011010";
            uut_rst <= '0';
          WHEN "00101011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101011011";
            uut_rst <= '0';
          WHEN "00101011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101011100";
            uut_rst <= '0';
          WHEN "00101011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101011101";
            uut_rst <= '0';
          WHEN "00101011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101011110";
            uut_rst <= '0';
          WHEN "00101011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101011111";
            uut_rst <= '0';
          WHEN "00101011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101100000";
            uut_rst <= '0';
          WHEN "00101100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101100001";
            uut_rst <= '0';
          WHEN "00101100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101100010";
            uut_rst <= '0';
          WHEN "00101100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101100011";
            uut_rst <= '0';
          WHEN "00101100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101100100";
            uut_rst <= '0';
          WHEN "00101100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101100101";
            uut_rst <= '0';
          WHEN "00101100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101100110";
            uut_rst <= '0';
          WHEN "00101100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101100111";
            uut_rst <= '0';
          WHEN "00101100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101101000";
            uut_rst <= '0';
          WHEN "00101101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101101001";
            uut_rst <= '0';
          WHEN "00101101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101101010";
            uut_rst <= '0';
          WHEN "00101101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101101011";
            uut_rst <= '0';
          WHEN "00101101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101101100";
            uut_rst <= '0';
          WHEN "00101101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101101101";
            uut_rst <= '0';
          WHEN "00101101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101101110";
            uut_rst <= '0';
          WHEN "00101101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101101111";
            uut_rst <= '0';
          WHEN "00101101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101110000";
            uut_rst <= '0';
          WHEN "00101110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101110001";
            uut_rst <= '0';
          WHEN "00101110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101110010";
            uut_rst <= '0';
          WHEN "00101110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101110011";
            uut_rst <= '0';
          WHEN "00101110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101110100";
            uut_rst <= '0';
          WHEN "00101110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101110101";
            uut_rst <= '0';
          WHEN "00101110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101110110";
            uut_rst <= '0';
          WHEN "00101110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101110111";
            uut_rst <= '0';
          WHEN "00101110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101111000";
            uut_rst <= '0';
          WHEN "00101111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101111001";
            uut_rst <= '0';
          WHEN "00101111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101111010";
            uut_rst <= '0';
          WHEN "00101111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101111011";
            uut_rst <= '0';
          WHEN "00101111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101111100";
            uut_rst <= '0';
          WHEN "00101111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101111101";
            uut_rst <= '0';
          WHEN "00101111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101111110";
            uut_rst <= '0';
          WHEN "00101111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00101111111";
            uut_rst <= '0';
          WHEN "00101111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110000000";
            uut_rst <= '0';
          WHEN "00110000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110000001";
            uut_rst <= '0';
          WHEN "00110000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110000010";
            uut_rst <= '0';
          WHEN "00110000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110000011";
            uut_rst <= '0';
          WHEN "00110000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110000100";
            uut_rst <= '0';
          WHEN "00110000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110000101";
            uut_rst <= '0';
          WHEN "00110000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110000110";
            uut_rst <= '0';
          WHEN "00110000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110000111";
            uut_rst <= '0';
          WHEN "00110000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110001000";
            uut_rst <= '0';
          WHEN "00110001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110001001";
            uut_rst <= '0';
          WHEN "00110001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110001010";
            uut_rst <= '0';
          WHEN "00110001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110001011";
            uut_rst <= '0';
          WHEN "00110001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110001100";
            uut_rst <= '0';
          WHEN "00110001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110001101";
            uut_rst <= '0';
          WHEN "00110001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110001110";
            uut_rst <= '0';
          WHEN "00110001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110001111";
            uut_rst <= '0';
          WHEN "00110001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110010000";
            uut_rst <= '0';
          WHEN "00110010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110010001";
            uut_rst <= '0';
          WHEN "00110010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110010010";
            uut_rst <= '0';
          WHEN "00110010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110010011";
            uut_rst <= '0';
          WHEN "00110010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110010100";
            uut_rst <= '0';
          WHEN "00110010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110010101";
            uut_rst <= '0';
          WHEN "00110010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110010110";
            uut_rst <= '0';
          WHEN "00110010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110010111";
            uut_rst <= '0';
          WHEN "00110010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110011000";
            uut_rst <= '0';
          WHEN "00110011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110011001";
            uut_rst <= '0';
          WHEN "00110011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110011010";
            uut_rst <= '0';
          WHEN "00110011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110011011";
            uut_rst <= '0';
          WHEN "00110011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110011100";
            uut_rst <= '0';
          WHEN "00110011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110011101";
            uut_rst <= '0';
          WHEN "00110011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110011110";
            uut_rst <= '0';
          WHEN "00110011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110011111";
            uut_rst <= '0';
          WHEN "00110011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110100000";
            uut_rst <= '0';
          WHEN "00110100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110100001";
            uut_rst <= '0';
          WHEN "00110100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110100010";
            uut_rst <= '0';
          WHEN "00110100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110100011";
            uut_rst <= '0';
          WHEN "00110100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110100100";
            uut_rst <= '0';
          WHEN "00110100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110100101";
            uut_rst <= '0';
          WHEN "00110100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110100110";
            uut_rst <= '0';
          WHEN "00110100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110100111";
            uut_rst <= '0';
          WHEN "00110100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110101000";
            uut_rst <= '0';
          WHEN "00110101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110101001";
            uut_rst <= '0';
          WHEN "00110101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110101010";
            uut_rst <= '0';
          WHEN "00110101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110101011";
            uut_rst <= '0';
          WHEN "00110101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110101100";
            uut_rst <= '0';
          WHEN "00110101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110101101";
            uut_rst <= '0';
          WHEN "00110101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110101110";
            uut_rst <= '0';
          WHEN "00110101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110101111";
            uut_rst <= '0';
          WHEN "00110101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110110000";
            uut_rst <= '0';
          WHEN "00110110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110110001";
            uut_rst <= '0';
          WHEN "00110110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110110010";
            uut_rst <= '0';
          WHEN "00110110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110110011";
            uut_rst <= '0';
          WHEN "00110110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110110100";
            uut_rst <= '0';
          WHEN "00110110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110110101";
            uut_rst <= '0';
          WHEN "00110110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110110110";
            uut_rst <= '0';
          WHEN "00110110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110110111";
            uut_rst <= '0';
          WHEN "00110110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110111000";
            uut_rst <= '0';
          WHEN "00110111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110111001";
            uut_rst <= '0';
          WHEN "00110111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110111010";
            uut_rst <= '0';
          WHEN "00110111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110111011";
            uut_rst <= '0';
          WHEN "00110111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110111100";
            uut_rst <= '0';
          WHEN "00110111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110111101";
            uut_rst <= '0';
          WHEN "00110111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110111110";
            uut_rst <= '0';
          WHEN "00110111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00110111111";
            uut_rst <= '0';
          WHEN "00110111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111000000";
            uut_rst <= '0';
          WHEN "00111000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111000001";
            uut_rst <= '0';
          WHEN "00111000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111000010";
            uut_rst <= '0';
          WHEN "00111000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111000011";
            uut_rst <= '0';
          WHEN "00111000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111000100";
            uut_rst <= '0';
          WHEN "00111000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111000101";
            uut_rst <= '0';
          WHEN "00111000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111000110";
            uut_rst <= '0';
          WHEN "00111000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111000111";
            uut_rst <= '0';
          WHEN "00111000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111001000";
            uut_rst <= '0';
          WHEN "00111001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111001001";
            uut_rst <= '0';
          WHEN "00111001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111001010";
            uut_rst <= '0';
          WHEN "00111001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111001011";
            uut_rst <= '0';
          WHEN "00111001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111001100";
            uut_rst <= '0';
          WHEN "00111001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111001101";
            uut_rst <= '0';
          WHEN "00111001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111001110";
            uut_rst <= '0';
          WHEN "00111001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111001111";
            uut_rst <= '0';
          WHEN "00111001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111010000";
            uut_rst <= '0';
          WHEN "00111010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111010001";
            uut_rst <= '0';
          WHEN "00111010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111010010";
            uut_rst <= '0';
          WHEN "00111010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111010011";
            uut_rst <= '0';
          WHEN "00111010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111010100";
            uut_rst <= '0';
          WHEN "00111010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111010101";
            uut_rst <= '0';
          WHEN "00111010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111010110";
            uut_rst <= '0';
          WHEN "00111010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111010111";
            uut_rst <= '0';
          WHEN "00111010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111011000";
            uut_rst <= '0';
          WHEN "00111011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111011001";
            uut_rst <= '0';
          WHEN "00111011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111011010";
            uut_rst <= '0';
          WHEN "00111011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111011011";
            uut_rst <= '0';
          WHEN "00111011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111011100";
            uut_rst <= '0';
          WHEN "00111011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111011101";
            uut_rst <= '0';
          WHEN "00111011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111011110";
            uut_rst <= '0';
          WHEN "00111011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111011111";
            uut_rst <= '0';
          WHEN "00111011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111100000";
            uut_rst <= '0';
          WHEN "00111100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111100001";
            uut_rst <= '0';
          WHEN "00111100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111100010";
            uut_rst <= '0';
          WHEN "00111100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111100011";
            uut_rst <= '0';
          WHEN "00111100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111100100";
            uut_rst <= '0';
          WHEN "00111100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111100101";
            uut_rst <= '0';
          WHEN "00111100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111100110";
            uut_rst <= '0';
          WHEN "00111100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111100111";
            uut_rst <= '0';
          WHEN "00111100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111101000";
            uut_rst <= '0';
          WHEN "00111101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111101001";
            uut_rst <= '0';
          WHEN "00111101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111101010";
            uut_rst <= '0';
          WHEN "00111101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111101011";
            uut_rst <= '0';
          WHEN "00111101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111101100";
            uut_rst <= '0';
          WHEN "00111101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111101101";
            uut_rst <= '0';
          WHEN "00111101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111101110";
            uut_rst <= '0';
          WHEN "00111101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111101111";
            uut_rst <= '0';
          WHEN "00111101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111110000";
            uut_rst <= '0';
          WHEN "00111110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111110001";
            uut_rst <= '0';
          WHEN "00111110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111110010";
            uut_rst <= '0';
          WHEN "00111110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111110011";
            uut_rst <= '0';
          WHEN "00111110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111110100";
            uut_rst <= '0';
          WHEN "00111110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111110101";
            uut_rst <= '0';
          WHEN "00111110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111110110";
            uut_rst <= '0';
          WHEN "00111110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111110111";
            uut_rst <= '0';
          WHEN "00111110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111111000";
            uut_rst <= '0';
          WHEN "00111111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111111001";
            uut_rst <= '0';
          WHEN "00111111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111111010";
            uut_rst <= '0';
          WHEN "00111111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111111011";
            uut_rst <= '0';
          WHEN "00111111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111111100";
            uut_rst <= '0';
          WHEN "00111111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111111101";
            uut_rst <= '0';
          WHEN "00111111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111111110";
            uut_rst <= '0';
          WHEN "00111111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "00111111111";
            uut_rst <= '0';
          WHEN "00111111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000000000";
            uut_rst <= '0';
          WHEN "01000000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000000001";
            uut_rst <= '0';
          WHEN "01000000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000000010";
            uut_rst <= '0';
          WHEN "01000000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000000011";
            uut_rst <= '0';
          WHEN "01000000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000000100";
            uut_rst <= '0';
          WHEN "01000000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000000101";
            uut_rst <= '0';
          WHEN "01000000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000000110";
            uut_rst <= '0';
          WHEN "01000000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000000111";
            uut_rst <= '0';
          WHEN "01000000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000001000";
            uut_rst <= '0';
          WHEN "01000001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000001001";
            uut_rst <= '0';
          WHEN "01000001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000001010";
            uut_rst <= '0';
          WHEN "01000001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000001011";
            uut_rst <= '0';
          WHEN "01000001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000001100";
            uut_rst <= '0';
          WHEN "01000001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000001101";
            uut_rst <= '0';
          WHEN "01000001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000001110";
            uut_rst <= '0';
          WHEN "01000001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000001111";
            uut_rst <= '0';
          WHEN "01000001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000010000";
            uut_rst <= '0';
          WHEN "01000010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000010001";
            uut_rst <= '0';
          WHEN "01000010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000010010";
            uut_rst <= '0';
          WHEN "01000010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000010011";
            uut_rst <= '0';
          WHEN "01000010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000010100";
            uut_rst <= '0';
          WHEN "01000010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000010101";
            uut_rst <= '0';
          WHEN "01000010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000010110";
            uut_rst <= '0';
          WHEN "01000010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000010111";
            uut_rst <= '0';
          WHEN "01000010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000011000";
            uut_rst <= '0';
          WHEN "01000011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000011001";
            uut_rst <= '0';
          WHEN "01000011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000011010";
            uut_rst <= '0';
          WHEN "01000011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000011011";
            uut_rst <= '0';
          WHEN "01000011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000011100";
            uut_rst <= '0';
          WHEN "01000011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000011101";
            uut_rst <= '0';
          WHEN "01000011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000011110";
            uut_rst <= '0';
          WHEN "01000011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000011111";
            uut_rst <= '0';
          WHEN "01000011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000100000";
            uut_rst <= '0';
          WHEN "01000100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000100001";
            uut_rst <= '0';
          WHEN "01000100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000100010";
            uut_rst <= '0';
          WHEN "01000100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000100011";
            uut_rst <= '0';
          WHEN "01000100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000100100";
            uut_rst <= '0';
          WHEN "01000100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000100101";
            uut_rst <= '0';
          WHEN "01000100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000100110";
            uut_rst <= '0';
          WHEN "01000100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000100111";
            uut_rst <= '0';
          WHEN "01000100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000101000";
            uut_rst <= '0';
          WHEN "01000101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000101001";
            uut_rst <= '0';
          WHEN "01000101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000101010";
            uut_rst <= '0';
          WHEN "01000101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000101011";
            uut_rst <= '0';
          WHEN "01000101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000101100";
            uut_rst <= '0';
          WHEN "01000101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000101101";
            uut_rst <= '0';
          WHEN "01000101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000101110";
            uut_rst <= '0';
          WHEN "01000101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000101111";
            uut_rst <= '0';
          WHEN "01000101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000110000";
            uut_rst <= '0';
          WHEN "01000110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000110001";
            uut_rst <= '0';
          WHEN "01000110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000110010";
            uut_rst <= '0';
          WHEN "01000110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000110011";
            uut_rst <= '0';
          WHEN "01000110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000110100";
            uut_rst <= '0';
          WHEN "01000110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000110101";
            uut_rst <= '0';
          WHEN "01000110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000110110";
            uut_rst <= '0';
          WHEN "01000110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000110111";
            uut_rst <= '0';
          WHEN "01000110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000111000";
            uut_rst <= '0';
          WHEN "01000111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000111001";
            uut_rst <= '0';
          WHEN "01000111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000111010";
            uut_rst <= '0';
          WHEN "01000111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000111011";
            uut_rst <= '0';
          WHEN "01000111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000111100";
            uut_rst <= '0';
          WHEN "01000111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000111101";
            uut_rst <= '0';
          WHEN "01000111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000111110";
            uut_rst <= '0';
          WHEN "01000111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01000111111";
            uut_rst <= '0';
          WHEN "01000111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001000000";
            uut_rst <= '0';
          WHEN "01001000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001000001";
            uut_rst <= '0';
          WHEN "01001000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001000010";
            uut_rst <= '0';
          WHEN "01001000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001000011";
            uut_rst <= '0';
          WHEN "01001000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001000100";
            uut_rst <= '0';
          WHEN "01001000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001000101";
            uut_rst <= '0';
          WHEN "01001000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001000110";
            uut_rst <= '0';
          WHEN "01001000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001000111";
            uut_rst <= '0';
          WHEN "01001000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001001000";
            uut_rst <= '0';
          WHEN "01001001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001001001";
            uut_rst <= '0';
          WHEN "01001001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001001010";
            uut_rst <= '0';
          WHEN "01001001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001001011";
            uut_rst <= '0';
          WHEN "01001001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001001100";
            uut_rst <= '0';
          WHEN "01001001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001001101";
            uut_rst <= '0';
          WHEN "01001001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001001110";
            uut_rst <= '0';
          WHEN "01001001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001001111";
            uut_rst <= '0';
          WHEN "01001001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001010000";
            uut_rst <= '0';
          WHEN "01001010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001010001";
            uut_rst <= '0';
          WHEN "01001010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001010010";
            uut_rst <= '0';
          WHEN "01001010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001010011";
            uut_rst <= '0';
          WHEN "01001010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001010100";
            uut_rst <= '0';
          WHEN "01001010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001010101";
            uut_rst <= '0';
          WHEN "01001010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001010110";
            uut_rst <= '0';
          WHEN "01001010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001010111";
            uut_rst <= '0';
          WHEN "01001010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001011000";
            uut_rst <= '0';
          WHEN "01001011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001011001";
            uut_rst <= '0';
          WHEN "01001011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001011010";
            uut_rst <= '0';
          WHEN "01001011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001011011";
            uut_rst <= '0';
          WHEN "01001011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001011100";
            uut_rst <= '0';
          WHEN "01001011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001011101";
            uut_rst <= '0';
          WHEN "01001011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001011110";
            uut_rst <= '0';
          WHEN "01001011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001011111";
            uut_rst <= '0';
          WHEN "01001011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001100000";
            uut_rst <= '0';
          WHEN "01001100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001100001";
            uut_rst <= '0';
          WHEN "01001100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001100010";
            uut_rst <= '0';
          WHEN "01001100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001100011";
            uut_rst <= '0';
          WHEN "01001100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001100100";
            uut_rst <= '0';
          WHEN "01001100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001100101";
            uut_rst <= '0';
          WHEN "01001100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001100110";
            uut_rst <= '0';
          WHEN "01001100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001100111";
            uut_rst <= '0';
          WHEN "01001100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001101000";
            uut_rst <= '0';
          WHEN "01001101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001101001";
            uut_rst <= '0';
          WHEN "01001101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001101010";
            uut_rst <= '0';
          WHEN "01001101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001101011";
            uut_rst <= '0';
          WHEN "01001101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001101100";
            uut_rst <= '0';
          WHEN "01001101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001101101";
            uut_rst <= '0';
          WHEN "01001101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001101110";
            uut_rst <= '0';
          WHEN "01001101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001101111";
            uut_rst <= '0';
          WHEN "01001101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001110000";
            uut_rst <= '0';
          WHEN "01001110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001110001";
            uut_rst <= '0';
          WHEN "01001110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001110010";
            uut_rst <= '0';
          WHEN "01001110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001110011";
            uut_rst <= '0';
          WHEN "01001110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001110100";
            uut_rst <= '0';
          WHEN "01001110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001110101";
            uut_rst <= '0';
          WHEN "01001110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001110110";
            uut_rst <= '0';
          WHEN "01001110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001110111";
            uut_rst <= '0';
          WHEN "01001110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001111000";
            uut_rst <= '0';
          WHEN "01001111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001111001";
            uut_rst <= '0';
          WHEN "01001111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001111010";
            uut_rst <= '0';
          WHEN "01001111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001111011";
            uut_rst <= '0';
          WHEN "01001111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001111100";
            uut_rst <= '0';
          WHEN "01001111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001111101";
            uut_rst <= '0';
          WHEN "01001111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001111110";
            uut_rst <= '0';
          WHEN "01001111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01001111111";
            uut_rst <= '0';
          WHEN "01001111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010000000";
            uut_rst <= '0';
          WHEN "01010000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010000001";
            uut_rst <= '0';
          WHEN "01010000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010000010";
            uut_rst <= '0';
          WHEN "01010000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010000011";
            uut_rst <= '0';
          WHEN "01010000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010000100";
            uut_rst <= '0';
          WHEN "01010000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010000101";
            uut_rst <= '0';
          WHEN "01010000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010000110";
            uut_rst <= '0';
          WHEN "01010000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010000111";
            uut_rst <= '0';
          WHEN "01010000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010001000";
            uut_rst <= '0';
          WHEN "01010001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010001001";
            uut_rst <= '0';
          WHEN "01010001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010001010";
            uut_rst <= '0';
          WHEN "01010001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010001011";
            uut_rst <= '0';
          WHEN "01010001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010001100";
            uut_rst <= '0';
          WHEN "01010001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010001101";
            uut_rst <= '0';
          WHEN "01010001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010001110";
            uut_rst <= '0';
          WHEN "01010001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010001111";
            uut_rst <= '0';
          WHEN "01010001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010010000";
            uut_rst <= '0';
          WHEN "01010010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010010001";
            uut_rst <= '0';
          WHEN "01010010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010010010";
            uut_rst <= '0';
          WHEN "01010010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010010011";
            uut_rst <= '0';
          WHEN "01010010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010010100";
            uut_rst <= '0';
          WHEN "01010010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010010101";
            uut_rst <= '0';
          WHEN "01010010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010010110";
            uut_rst <= '0';
          WHEN "01010010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010010111";
            uut_rst <= '0';
          WHEN "01010010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010011000";
            uut_rst <= '0';
          WHEN "01010011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010011001";
            uut_rst <= '0';
          WHEN "01010011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010011010";
            uut_rst <= '0';
          WHEN "01010011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010011011";
            uut_rst <= '0';
          WHEN "01010011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010011100";
            uut_rst <= '0';
          WHEN "01010011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010011101";
            uut_rst <= '0';
          WHEN "01010011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010011110";
            uut_rst <= '0';
          WHEN "01010011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010011111";
            uut_rst <= '0';
          WHEN "01010011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010100000";
            uut_rst <= '0';
          WHEN "01010100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010100001";
            uut_rst <= '0';
          WHEN "01010100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010100010";
            uut_rst <= '0';
          WHEN "01010100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010100011";
            uut_rst <= '0';
          WHEN "01010100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010100100";
            uut_rst <= '0';
          WHEN "01010100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010100101";
            uut_rst <= '0';
          WHEN "01010100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010100110";
            uut_rst <= '0';
          WHEN "01010100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010100111";
            uut_rst <= '0';
          WHEN "01010100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010101000";
            uut_rst <= '0';
          WHEN "01010101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010101001";
            uut_rst <= '0';
          WHEN "01010101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010101010";
            uut_rst <= '0';
          WHEN "01010101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010101011";
            uut_rst <= '0';
          WHEN "01010101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010101100";
            uut_rst <= '0';
          WHEN "01010101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010101101";
            uut_rst <= '0';
          WHEN "01010101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010101110";
            uut_rst <= '0';
          WHEN "01010101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010101111";
            uut_rst <= '0';
          WHEN "01010101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010110000";
            uut_rst <= '0';
          WHEN "01010110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010110001";
            uut_rst <= '0';
          WHEN "01010110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010110010";
            uut_rst <= '0';
          WHEN "01010110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010110011";
            uut_rst <= '0';
          WHEN "01010110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010110100";
            uut_rst <= '0';
          WHEN "01010110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010110101";
            uut_rst <= '0';
          WHEN "01010110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010110110";
            uut_rst <= '0';
          WHEN "01010110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010110111";
            uut_rst <= '0';
          WHEN "01010110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010111000";
            uut_rst <= '0';
          WHEN "01010111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010111001";
            uut_rst <= '0';
          WHEN "01010111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010111010";
            uut_rst <= '0';
          WHEN "01010111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010111011";
            uut_rst <= '0';
          WHEN "01010111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010111100";
            uut_rst <= '0';
          WHEN "01010111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010111101";
            uut_rst <= '0';
          WHEN "01010111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010111110";
            uut_rst <= '0';
          WHEN "01010111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01010111111";
            uut_rst <= '0';
          WHEN "01010111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011000000";
            uut_rst <= '0';
          WHEN "01011000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011000001";
            uut_rst <= '0';
          WHEN "01011000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011000010";
            uut_rst <= '0';
          WHEN "01011000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011000011";
            uut_rst <= '0';
          WHEN "01011000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011000100";
            uut_rst <= '0';
          WHEN "01011000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011000101";
            uut_rst <= '0';
          WHEN "01011000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011000110";
            uut_rst <= '0';
          WHEN "01011000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011000111";
            uut_rst <= '0';
          WHEN "01011000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011001000";
            uut_rst <= '0';
          WHEN "01011001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011001001";
            uut_rst <= '0';
          WHEN "01011001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011001010";
            uut_rst <= '0';
          WHEN "01011001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011001011";
            uut_rst <= '0';
          WHEN "01011001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011001100";
            uut_rst <= '0';
          WHEN "01011001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011001101";
            uut_rst <= '0';
          WHEN "01011001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011001110";
            uut_rst <= '0';
          WHEN "01011001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011001111";
            uut_rst <= '0';
          WHEN "01011001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011010000";
            uut_rst <= '0';
          WHEN "01011010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011010001";
            uut_rst <= '0';
          WHEN "01011010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011010010";
            uut_rst <= '0';
          WHEN "01011010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011010011";
            uut_rst <= '0';
          WHEN "01011010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011010100";
            uut_rst <= '0';
          WHEN "01011010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011010101";
            uut_rst <= '0';
          WHEN "01011010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011010110";
            uut_rst <= '0';
          WHEN "01011010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011010111";
            uut_rst <= '0';
          WHEN "01011010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011011000";
            uut_rst <= '0';
          WHEN "01011011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011011001";
            uut_rst <= '0';
          WHEN "01011011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011011010";
            uut_rst <= '0';
          WHEN "01011011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011011011";
            uut_rst <= '0';
          WHEN "01011011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011011100";
            uut_rst <= '0';
          WHEN "01011011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011011101";
            uut_rst <= '0';
          WHEN "01011011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011011110";
            uut_rst <= '0';
          WHEN "01011011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011011111";
            uut_rst <= '0';
          WHEN "01011011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011100000";
            uut_rst <= '0';
          WHEN "01011100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011100001";
            uut_rst <= '0';
          WHEN "01011100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011100010";
            uut_rst <= '0';
          WHEN "01011100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011100011";
            uut_rst <= '0';
          WHEN "01011100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011100100";
            uut_rst <= '0';
          WHEN "01011100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011100101";
            uut_rst <= '0';
          WHEN "01011100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011100110";
            uut_rst <= '0';
          WHEN "01011100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011100111";
            uut_rst <= '0';
          WHEN "01011100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011101000";
            uut_rst <= '0';
          WHEN "01011101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011101001";
            uut_rst <= '0';
          WHEN "01011101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011101010";
            uut_rst <= '0';
          WHEN "01011101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011101011";
            uut_rst <= '0';
          WHEN "01011101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011101100";
            uut_rst <= '0';
          WHEN "01011101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011101101";
            uut_rst <= '0';
          WHEN "01011101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011101110";
            uut_rst <= '0';
          WHEN "01011101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011101111";
            uut_rst <= '0';
          WHEN "01011101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011110000";
            uut_rst <= '0';
          WHEN "01011110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011110001";
            uut_rst <= '0';
          WHEN "01011110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011110010";
            uut_rst <= '0';
          WHEN "01011110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011110011";
            uut_rst <= '0';
          WHEN "01011110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011110100";
            uut_rst <= '0';
          WHEN "01011110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011110101";
            uut_rst <= '0';
          WHEN "01011110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011110110";
            uut_rst <= '0';
          WHEN "01011110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011110111";
            uut_rst <= '0';
          WHEN "01011110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011111000";
            uut_rst <= '0';
          WHEN "01011111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011111001";
            uut_rst <= '0';
          WHEN "01011111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011111010";
            uut_rst <= '0';
          WHEN "01011111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011111011";
            uut_rst <= '0';
          WHEN "01011111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011111100";
            uut_rst <= '0';
          WHEN "01011111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011111101";
            uut_rst <= '0';
          WHEN "01011111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011111110";
            uut_rst <= '0';
          WHEN "01011111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01011111111";
            uut_rst <= '0';
          WHEN "01011111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100000000";
            uut_rst <= '0';
          WHEN "01100000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100000001";
            uut_rst <= '0';
          WHEN "01100000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100000010";
            uut_rst <= '0';
          WHEN "01100000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100000011";
            uut_rst <= '0';
          WHEN "01100000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100000100";
            uut_rst <= '0';
          WHEN "01100000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100000101";
            uut_rst <= '0';
          WHEN "01100000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100000110";
            uut_rst <= '0';
          WHEN "01100000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100000111";
            uut_rst <= '0';
          WHEN "01100000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100001000";
            uut_rst <= '0';
          WHEN "01100001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100001001";
            uut_rst <= '0';
          WHEN "01100001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100001010";
            uut_rst <= '0';
          WHEN "01100001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100001011";
            uut_rst <= '0';
          WHEN "01100001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100001100";
            uut_rst <= '0';
          WHEN "01100001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100001101";
            uut_rst <= '0';
          WHEN "01100001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100001110";
            uut_rst <= '0';
          WHEN "01100001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100001111";
            uut_rst <= '0';
          WHEN "01100001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100010000";
            uut_rst <= '0';
          WHEN "01100010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100010001";
            uut_rst <= '0';
          WHEN "01100010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100010010";
            uut_rst <= '0';
          WHEN "01100010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100010011";
            uut_rst <= '0';
          WHEN "01100010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100010100";
            uut_rst <= '0';
          WHEN "01100010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100010101";
            uut_rst <= '0';
          WHEN "01100010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100010110";
            uut_rst <= '0';
          WHEN "01100010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100010111";
            uut_rst <= '0';
          WHEN "01100010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100011000";
            uut_rst <= '0';
          WHEN "01100011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100011001";
            uut_rst <= '0';
          WHEN "01100011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100011010";
            uut_rst <= '0';
          WHEN "01100011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100011011";
            uut_rst <= '0';
          WHEN "01100011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100011100";
            uut_rst <= '0';
          WHEN "01100011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100011101";
            uut_rst <= '0';
          WHEN "01100011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100011110";
            uut_rst <= '0';
          WHEN "01100011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100011111";
            uut_rst <= '0';
          WHEN "01100011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100100000";
            uut_rst <= '0';
          WHEN "01100100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100100001";
            uut_rst <= '0';
          WHEN "01100100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100100010";
            uut_rst <= '0';
          WHEN "01100100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100100011";
            uut_rst <= '0';
          WHEN "01100100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100100100";
            uut_rst <= '0';
          WHEN "01100100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100100101";
            uut_rst <= '0';
          WHEN "01100100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100100110";
            uut_rst <= '0';
          WHEN "01100100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100100111";
            uut_rst <= '0';
          WHEN "01100100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100101000";
            uut_rst <= '0';
          WHEN "01100101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100101001";
            uut_rst <= '0';
          WHEN "01100101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100101010";
            uut_rst <= '0';
          WHEN "01100101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100101011";
            uut_rst <= '0';
          WHEN "01100101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100101100";
            uut_rst <= '0';
          WHEN "01100101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100101101";
            uut_rst <= '0';
          WHEN "01100101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100101110";
            uut_rst <= '0';
          WHEN "01100101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100101111";
            uut_rst <= '0';
          WHEN "01100101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100110000";
            uut_rst <= '0';
          WHEN "01100110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100110001";
            uut_rst <= '0';
          WHEN "01100110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100110010";
            uut_rst <= '0';
          WHEN "01100110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100110011";
            uut_rst <= '0';
          WHEN "01100110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100110100";
            uut_rst <= '0';
          WHEN "01100110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100110101";
            uut_rst <= '0';
          WHEN "01100110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100110110";
            uut_rst <= '0';
          WHEN "01100110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100110111";
            uut_rst <= '0';
          WHEN "01100110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100111000";
            uut_rst <= '0';
          WHEN "01100111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100111001";
            uut_rst <= '0';
          WHEN "01100111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100111010";
            uut_rst <= '0';
          WHEN "01100111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100111011";
            uut_rst <= '0';
          WHEN "01100111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100111100";
            uut_rst <= '0';
          WHEN "01100111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100111101";
            uut_rst <= '0';
          WHEN "01100111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100111110";
            uut_rst <= '0';
          WHEN "01100111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01100111111";
            uut_rst <= '0';
          WHEN "01100111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101000000";
            uut_rst <= '0';
          WHEN "01101000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101000001";
            uut_rst <= '0';
          WHEN "01101000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101000010";
            uut_rst <= '0';
          WHEN "01101000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101000011";
            uut_rst <= '0';
          WHEN "01101000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101000100";
            uut_rst <= '0';
          WHEN "01101000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101000101";
            uut_rst <= '0';
          WHEN "01101000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101000110";
            uut_rst <= '0';
          WHEN "01101000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101000111";
            uut_rst <= '0';
          WHEN "01101000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101001000";
            uut_rst <= '0';
          WHEN "01101001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101001001";
            uut_rst <= '0';
          WHEN "01101001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101001010";
            uut_rst <= '0';
          WHEN "01101001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101001011";
            uut_rst <= '0';
          WHEN "01101001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101001100";
            uut_rst <= '0';
          WHEN "01101001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101001101";
            uut_rst <= '0';
          WHEN "01101001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101001110";
            uut_rst <= '0';
          WHEN "01101001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101001111";
            uut_rst <= '0';
          WHEN "01101001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101010000";
            uut_rst <= '0';
          WHEN "01101010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101010001";
            uut_rst <= '0';
          WHEN "01101010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101010010";
            uut_rst <= '0';
          WHEN "01101010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101010011";
            uut_rst <= '0';
          WHEN "01101010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101010100";
            uut_rst <= '0';
          WHEN "01101010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101010101";
            uut_rst <= '0';
          WHEN "01101010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101010110";
            uut_rst <= '0';
          WHEN "01101010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101010111";
            uut_rst <= '0';
          WHEN "01101010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101011000";
            uut_rst <= '0';
          WHEN "01101011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101011001";
            uut_rst <= '0';
          WHEN "01101011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101011010";
            uut_rst <= '0';
          WHEN "01101011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101011011";
            uut_rst <= '0';
          WHEN "01101011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101011100";
            uut_rst <= '0';
          WHEN "01101011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101011101";
            uut_rst <= '0';
          WHEN "01101011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101011110";
            uut_rst <= '0';
          WHEN "01101011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101011111";
            uut_rst <= '0';
          WHEN "01101011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101100000";
            uut_rst <= '0';
          WHEN "01101100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101100001";
            uut_rst <= '0';
          WHEN "01101100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101100010";
            uut_rst <= '0';
          WHEN "01101100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101100011";
            uut_rst <= '0';
          WHEN "01101100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101100100";
            uut_rst <= '0';
          WHEN "01101100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101100101";
            uut_rst <= '0';
          WHEN "01101100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101100110";
            uut_rst <= '0';
          WHEN "01101100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101100111";
            uut_rst <= '0';
          WHEN "01101100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101101000";
            uut_rst <= '0';
          WHEN "01101101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101101001";
            uut_rst <= '0';
          WHEN "01101101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101101010";
            uut_rst <= '0';
          WHEN "01101101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101101011";
            uut_rst <= '0';
          WHEN "01101101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101101100";
            uut_rst <= '0';
          WHEN "01101101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101101101";
            uut_rst <= '0';
          WHEN "01101101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101101110";
            uut_rst <= '0';
          WHEN "01101101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101101111";
            uut_rst <= '0';
          WHEN "01101101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101110000";
            uut_rst <= '0';
          WHEN "01101110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101110001";
            uut_rst <= '0';
          WHEN "01101110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101110010";
            uut_rst <= '0';
          WHEN "01101110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101110011";
            uut_rst <= '0';
          WHEN "01101110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101110100";
            uut_rst <= '0';
          WHEN "01101110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101110101";
            uut_rst <= '0';
          WHEN "01101110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101110110";
            uut_rst <= '0';
          WHEN "01101110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101110111";
            uut_rst <= '0';
          WHEN "01101110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101111000";
            uut_rst <= '0';
          WHEN "01101111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101111001";
            uut_rst <= '0';
          WHEN "01101111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101111010";
            uut_rst <= '0';
          WHEN "01101111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101111011";
            uut_rst <= '0';
          WHEN "01101111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101111100";
            uut_rst <= '0';
          WHEN "01101111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101111101";
            uut_rst <= '0';
          WHEN "01101111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101111110";
            uut_rst <= '0';
          WHEN "01101111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01101111111";
            uut_rst <= '0';
          WHEN "01101111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110000000";
            uut_rst <= '0';
          WHEN "01110000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110000001";
            uut_rst <= '0';
          WHEN "01110000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110000010";
            uut_rst <= '0';
          WHEN "01110000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110000011";
            uut_rst <= '0';
          WHEN "01110000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110000100";
            uut_rst <= '0';
          WHEN "01110000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110000101";
            uut_rst <= '0';
          WHEN "01110000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110000110";
            uut_rst <= '0';
          WHEN "01110000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110000111";
            uut_rst <= '0';
          WHEN "01110000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110001000";
            uut_rst <= '0';
          WHEN "01110001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110001001";
            uut_rst <= '0';
          WHEN "01110001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110001010";
            uut_rst <= '0';
          WHEN "01110001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110001011";
            uut_rst <= '0';
          WHEN "01110001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110001100";
            uut_rst <= '0';
          WHEN "01110001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110001101";
            uut_rst <= '0';
          WHEN "01110001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110001110";
            uut_rst <= '0';
          WHEN "01110001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110001111";
            uut_rst <= '0';
          WHEN "01110001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110010000";
            uut_rst <= '0';
          WHEN "01110010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110010001";
            uut_rst <= '0';
          WHEN "01110010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110010010";
            uut_rst <= '0';
          WHEN "01110010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110010011";
            uut_rst <= '0';
          WHEN "01110010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110010100";
            uut_rst <= '0';
          WHEN "01110010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110010101";
            uut_rst <= '0';
          WHEN "01110010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110010110";
            uut_rst <= '0';
          WHEN "01110010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110010111";
            uut_rst <= '0';
          WHEN "01110010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110011000";
            uut_rst <= '0';
          WHEN "01110011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110011001";
            uut_rst <= '0';
          WHEN "01110011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110011010";
            uut_rst <= '0';
          WHEN "01110011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110011011";
            uut_rst <= '0';
          WHEN "01110011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110011100";
            uut_rst <= '0';
          WHEN "01110011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110011101";
            uut_rst <= '0';
          WHEN "01110011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110011110";
            uut_rst <= '0';
          WHEN "01110011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110011111";
            uut_rst <= '0';
          WHEN "01110011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110100000";
            uut_rst <= '0';
          WHEN "01110100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110100001";
            uut_rst <= '0';
          WHEN "01110100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110100010";
            uut_rst <= '0';
          WHEN "01110100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110100011";
            uut_rst <= '0';
          WHEN "01110100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110100100";
            uut_rst <= '0';
          WHEN "01110100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110100101";
            uut_rst <= '0';
          WHEN "01110100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110100110";
            uut_rst <= '0';
          WHEN "01110100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110100111";
            uut_rst <= '0';
          WHEN "01110100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110101000";
            uut_rst <= '0';
          WHEN "01110101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110101001";
            uut_rst <= '0';
          WHEN "01110101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110101010";
            uut_rst <= '0';
          WHEN "01110101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110101011";
            uut_rst <= '0';
          WHEN "01110101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110101100";
            uut_rst <= '0';
          WHEN "01110101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110101101";
            uut_rst <= '0';
          WHEN "01110101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110101110";
            uut_rst <= '0';
          WHEN "01110101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110101111";
            uut_rst <= '0';
          WHEN "01110101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110110000";
            uut_rst <= '0';
          WHEN "01110110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110110001";
            uut_rst <= '0';
          WHEN "01110110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110110010";
            uut_rst <= '0';
          WHEN "01110110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110110011";
            uut_rst <= '0';
          WHEN "01110110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110110100";
            uut_rst <= '0';
          WHEN "01110110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110110101";
            uut_rst <= '0';
          WHEN "01110110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110110110";
            uut_rst <= '0';
          WHEN "01110110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110110111";
            uut_rst <= '0';
          WHEN "01110110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110111000";
            uut_rst <= '0';
          WHEN "01110111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110111001";
            uut_rst <= '0';
          WHEN "01110111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110111010";
            uut_rst <= '0';
          WHEN "01110111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110111011";
            uut_rst <= '0';
          WHEN "01110111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110111100";
            uut_rst <= '0';
          WHEN "01110111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110111101";
            uut_rst <= '0';
          WHEN "01110111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110111110";
            uut_rst <= '0';
          WHEN "01110111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01110111111";
            uut_rst <= '0';
          WHEN "01110111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111000000";
            uut_rst <= '0';
          WHEN "01111000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111000001";
            uut_rst <= '0';
          WHEN "01111000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111000010";
            uut_rst <= '0';
          WHEN "01111000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111000011";
            uut_rst <= '0';
          WHEN "01111000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111000100";
            uut_rst <= '0';
          WHEN "01111000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111000101";
            uut_rst <= '0';
          WHEN "01111000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111000110";
            uut_rst <= '0';
          WHEN "01111000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111000111";
            uut_rst <= '0';
          WHEN "01111000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111001000";
            uut_rst <= '0';
          WHEN "01111001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111001001";
            uut_rst <= '0';
          WHEN "01111001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111001010";
            uut_rst <= '0';
          WHEN "01111001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111001011";
            uut_rst <= '0';
          WHEN "01111001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111001100";
            uut_rst <= '0';
          WHEN "01111001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111001101";
            uut_rst <= '0';
          WHEN "01111001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111001110";
            uut_rst <= '0';
          WHEN "01111001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111001111";
            uut_rst <= '0';
          WHEN "01111001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111010000";
            uut_rst <= '0';
          WHEN "01111010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111010001";
            uut_rst <= '0';
          WHEN "01111010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111010010";
            uut_rst <= '0';
          WHEN "01111010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111010011";
            uut_rst <= '0';
          WHEN "01111010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111010100";
            uut_rst <= '0';
          WHEN "01111010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111010101";
            uut_rst <= '0';
          WHEN "01111010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111010110";
            uut_rst <= '0';
          WHEN "01111010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111010111";
            uut_rst <= '0';
          WHEN "01111010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111011000";
            uut_rst <= '0';
          WHEN "01111011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111011001";
            uut_rst <= '0';
          WHEN "01111011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111011010";
            uut_rst <= '0';
          WHEN "01111011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111011011";
            uut_rst <= '0';
          WHEN "01111011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111011100";
            uut_rst <= '0';
          WHEN "01111011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111011101";
            uut_rst <= '0';
          WHEN "01111011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111011110";
            uut_rst <= '0';
          WHEN "01111011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111011111";
            uut_rst <= '0';
          WHEN "01111011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111100000";
            uut_rst <= '0';
          WHEN "01111100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111100001";
            uut_rst <= '0';
          WHEN "01111100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111100010";
            uut_rst <= '0';
          WHEN "01111100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111100011";
            uut_rst <= '0';
          WHEN "01111100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111100100";
            uut_rst <= '0';
          WHEN "01111100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111100101";
            uut_rst <= '0';
          WHEN "01111100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111100110";
            uut_rst <= '0';
          WHEN "01111100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111100111";
            uut_rst <= '0';
          WHEN "01111100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111101000";
            uut_rst <= '0';
          WHEN "01111101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111101001";
            uut_rst <= '0';
          WHEN "01111101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111101010";
            uut_rst <= '0';
          WHEN "01111101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111101011";
            uut_rst <= '0';
          WHEN "01111101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111101100";
            uut_rst <= '0';
          WHEN "01111101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111101101";
            uut_rst <= '0';
          WHEN "01111101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111101110";
            uut_rst <= '0';
          WHEN "01111101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111101111";
            uut_rst <= '0';
          WHEN "01111101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111110000";
            uut_rst <= '0';
          WHEN "01111110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111110001";
            uut_rst <= '0';
          WHEN "01111110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111110010";
            uut_rst <= '0';
          WHEN "01111110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111110011";
            uut_rst <= '0';
          WHEN "01111110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111110100";
            uut_rst <= '0';
          WHEN "01111110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111110101";
            uut_rst <= '0';
          WHEN "01111110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111110110";
            uut_rst <= '0';
          WHEN "01111110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111110111";
            uut_rst <= '0';
          WHEN "01111110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111111000";
            uut_rst <= '0';
          WHEN "01111111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111111001";
            uut_rst <= '0';
          WHEN "01111111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111111010";
            uut_rst <= '0';
          WHEN "01111111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111111011";
            uut_rst <= '0';
          WHEN "01111111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111111100";
            uut_rst <= '0';
          WHEN "01111111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111111101";
            uut_rst <= '0';
          WHEN "01111111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111111110";
            uut_rst <= '0';
          WHEN "01111111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "01111111111";
            uut_rst <= '0';
          WHEN "01111111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000000000";
            uut_rst <= '0';
          WHEN "10000000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000000001";
            uut_rst <= '0';
          WHEN "10000000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000000010";
            uut_rst <= '0';
          WHEN "10000000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000000011";
            uut_rst <= '0';
          WHEN "10000000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000000100";
            uut_rst <= '0';
          WHEN "10000000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000000101";
            uut_rst <= '0';
          WHEN "10000000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000000110";
            uut_rst <= '0';
          WHEN "10000000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000000111";
            uut_rst <= '0';
          WHEN "10000000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000001000";
            uut_rst <= '0';
          WHEN "10000001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000001001";
            uut_rst <= '0';
          WHEN "10000001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000001010";
            uut_rst <= '0';
          WHEN "10000001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000001011";
            uut_rst <= '0';
          WHEN "10000001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000001100";
            uut_rst <= '0';
          WHEN "10000001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000001101";
            uut_rst <= '0';
          WHEN "10000001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000001110";
            uut_rst <= '0';
          WHEN "10000001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000001111";
            uut_rst <= '0';
          WHEN "10000001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000010000";
            uut_rst <= '0';
          WHEN "10000010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000010001";
            uut_rst <= '0';
          WHEN "10000010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000010010";
            uut_rst <= '0';
          WHEN "10000010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000010011";
            uut_rst <= '0';
          WHEN "10000010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000010100";
            uut_rst <= '0';
          WHEN "10000010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000010101";
            uut_rst <= '0';
          WHEN "10000010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000010110";
            uut_rst <= '0';
          WHEN "10000010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000010111";
            uut_rst <= '0';
          WHEN "10000010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000011000";
            uut_rst <= '0';
          WHEN "10000011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000011001";
            uut_rst <= '0';
          WHEN "10000011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000011010";
            uut_rst <= '0';
          WHEN "10000011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000011011";
            uut_rst <= '0';
          WHEN "10000011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000011100";
            uut_rst <= '0';
          WHEN "10000011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000011101";
            uut_rst <= '0';
          WHEN "10000011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000011110";
            uut_rst <= '0';
          WHEN "10000011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000011111";
            uut_rst <= '0';
          WHEN "10000011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000100000";
            uut_rst <= '0';
          WHEN "10000100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000100001";
            uut_rst <= '0';
          WHEN "10000100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000100010";
            uut_rst <= '0';
          WHEN "10000100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000100011";
            uut_rst <= '0';
          WHEN "10000100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000100100";
            uut_rst <= '0';
          WHEN "10000100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000100101";
            uut_rst <= '0';
          WHEN "10000100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000100110";
            uut_rst <= '0';
          WHEN "10000100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000100111";
            uut_rst <= '0';
          WHEN "10000100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000101000";
            uut_rst <= '0';
          WHEN "10000101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000101001";
            uut_rst <= '0';
          WHEN "10000101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000101010";
            uut_rst <= '0';
          WHEN "10000101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000101011";
            uut_rst <= '0';
          WHEN "10000101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000101100";
            uut_rst <= '0';
          WHEN "10000101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000101101";
            uut_rst <= '0';
          WHEN "10000101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000101110";
            uut_rst <= '0';
          WHEN "10000101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000101111";
            uut_rst <= '0';
          WHEN "10000101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000110000";
            uut_rst <= '0';
          WHEN "10000110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000110001";
            uut_rst <= '0';
          WHEN "10000110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000110010";
            uut_rst <= '0';
          WHEN "10000110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000110011";
            uut_rst <= '0';
          WHEN "10000110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000110100";
            uut_rst <= '0';
          WHEN "10000110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000110101";
            uut_rst <= '0';
          WHEN "10000110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000110110";
            uut_rst <= '0';
          WHEN "10000110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000110111";
            uut_rst <= '0';
          WHEN "10000110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000111000";
            uut_rst <= '0';
          WHEN "10000111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000111001";
            uut_rst <= '0';
          WHEN "10000111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000111010";
            uut_rst <= '0';
          WHEN "10000111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000111011";
            uut_rst <= '0';
          WHEN "10000111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000111100";
            uut_rst <= '0';
          WHEN "10000111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000111101";
            uut_rst <= '0';
          WHEN "10000111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000111110";
            uut_rst <= '0';
          WHEN "10000111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10000111111";
            uut_rst <= '0';
          WHEN "10000111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001000000";
            uut_rst <= '0';
          WHEN "10001000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001000001";
            uut_rst <= '0';
          WHEN "10001000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001000010";
            uut_rst <= '0';
          WHEN "10001000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001000011";
            uut_rst <= '0';
          WHEN "10001000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001000100";
            uut_rst <= '0';
          WHEN "10001000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001000101";
            uut_rst <= '0';
          WHEN "10001000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001000110";
            uut_rst <= '0';
          WHEN "10001000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001000111";
            uut_rst <= '0';
          WHEN "10001000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001001000";
            uut_rst <= '0';
          WHEN "10001001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001001001";
            uut_rst <= '0';
          WHEN "10001001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001001010";
            uut_rst <= '0';
          WHEN "10001001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001001011";
            uut_rst <= '0';
          WHEN "10001001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001001100";
            uut_rst <= '0';
          WHEN "10001001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001001101";
            uut_rst <= '0';
          WHEN "10001001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001001110";
            uut_rst <= '0';
          WHEN "10001001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001001111";
            uut_rst <= '0';
          WHEN "10001001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001010000";
            uut_rst <= '0';
          WHEN "10001010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001010001";
            uut_rst <= '0';
          WHEN "10001010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001010010";
            uut_rst <= '0';
          WHEN "10001010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001010011";
            uut_rst <= '0';
          WHEN "10001010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001010100";
            uut_rst <= '0';
          WHEN "10001010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001010101";
            uut_rst <= '0';
          WHEN "10001010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001010110";
            uut_rst <= '0';
          WHEN "10001010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001010111";
            uut_rst <= '0';
          WHEN "10001010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001011000";
            uut_rst <= '0';
          WHEN "10001011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001011001";
            uut_rst <= '0';
          WHEN "10001011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001011010";
            uut_rst <= '0';
          WHEN "10001011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001011011";
            uut_rst <= '0';
          WHEN "10001011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001011100";
            uut_rst <= '0';
          WHEN "10001011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001011101";
            uut_rst <= '0';
          WHEN "10001011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001011110";
            uut_rst <= '0';
          WHEN "10001011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001011111";
            uut_rst <= '0';
          WHEN "10001011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001100000";
            uut_rst <= '0';
          WHEN "10001100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001100001";
            uut_rst <= '0';
          WHEN "10001100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001100010";
            uut_rst <= '0';
          WHEN "10001100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001100011";
            uut_rst <= '0';
          WHEN "10001100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001100100";
            uut_rst <= '0';
          WHEN "10001100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001100101";
            uut_rst <= '0';
          WHEN "10001100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001100110";
            uut_rst <= '0';
          WHEN "10001100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001100111";
            uut_rst <= '0';
          WHEN "10001100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001101000";
            uut_rst <= '0';
          WHEN "10001101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001101001";
            uut_rst <= '0';
          WHEN "10001101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001101010";
            uut_rst <= '0';
          WHEN "10001101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001101011";
            uut_rst <= '0';
          WHEN "10001101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001101100";
            uut_rst <= '0';
          WHEN "10001101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "10001101101";
            uut_rst <= '0';
          WHEN "10001101101" =>
            state <= "10001101110";
            uut_rst <= '0';
          WHEN "10001101110" =>
            state <= "10001101111";
            uut_rst <= '0';
          WHEN "10001101111" =>
            state <= "10001110000";
            uut_rst <= '0';
          WHEN "10001110000" =>
            state <= "10001110001";
            uut_rst <= '0';
          WHEN "10001110001" =>
            state <= "10001110010";
            uut_rst <= '0';
          WHEN "10001110010" =>
            state <= "10001110011";
            uut_rst <= '0';
          WHEN "10001110011" =>
            state <= "10001110100";
            uut_rst <= '0';
          WHEN "10001110100" =>
            state <= "10001110101";
            uut_rst <= '0';
          WHEN "10001110101" =>
            state <= "10001110110";
            uut_rst <= '0';
          WHEN "10001110110" =>
            state <= "10001110111";
            uut_rst <= '0';
          WHEN "10001110111" =>
            state <= "10001111000";
            uut_rst <= '0';
          WHEN "10001111000" =>
            state <= "10001111001";
            uut_rst <= '0';
          WHEN "10001111001" =>
            state <= "10001111010";
            uut_rst <= '0';
          WHEN "10001111010" =>
            state <= "10001111011";
            uut_rst <= '0';
          WHEN "10001111011" =>
            state <= "10001111100";
            uut_rst <= '0';
          WHEN "10001111100" =>
            state <= "10001111101";
            uut_rst <= '0';
          WHEN "10001111101" =>
            state <= "10001111110";
            uut_rst <= '0';
          WHEN "10001111110" =>
            state <= "10001111111";
            uut_rst <= '0';
          WHEN "10001111111" =>
            state <= "10010000000";
            uut_rst <= '0';
          WHEN "10010000000" =>
            state <= "10010000001";
            uut_rst <= '0';
          WHEN "10010000001" =>
            state <= "10010000010";
            uut_rst <= '0';
          WHEN "10010000010" =>
            state <= "10010000011";
            uut_rst <= '0';
          WHEN "10010000011" =>
            state <= "10010000100";
            uut_rst <= '0';
          WHEN "10010000100" =>
            state <= "10010000101";
            uut_rst <= '0';
          WHEN "10010000101" =>
            state <= "10010000110";
            uut_rst <= '0';
          WHEN "10010000110" =>
            state <= "10010000111";
            uut_rst <= '0';
          WHEN "10010000111" =>
            state <= "10010001000";
            uut_rst <= '0';
          WHEN "10010001000" =>
            state <= "10010001001";
            uut_rst <= '0';
          WHEN "10010001001" =>
            state <= "10010001010";
            uut_rst <= '0';
          WHEN "10010001010" =>
            state <= "10010001011";
            uut_rst <= '0';
          WHEN "10010001011" =>
            state <= "10010001100";
            uut_rst <= '0';
          WHEN "10010001100" =>
            state <= "10010001101";
            uut_rst <= '0';
          WHEN "10010001101" =>
            state <= "10010001110";
            uut_rst <= '0';
          WHEN "10010001110" =>
            state <= "10010001111";
            uut_rst <= '0';
          WHEN "10010001111" =>
            state <= "10010010000";
            uut_rst <= '0';
          WHEN "10010010000" =>
            state <= "10010010001";
            uut_rst <= '0';
          WHEN "10010010001" =>
            state <= "10010010010";
            uut_rst <= '0';
          WHEN "10010010010" =>
            state <= "10010010011";
            uut_rst <= '0';
          WHEN "10010010011" =>
            state <= "10010010100";
            uut_rst <= '0';
          WHEN "10010010100" =>
            state <= "10010010101";
            uut_rst <= '0';
          WHEN "10010010101" =>
            state <= "10010010110";
            uut_rst <= '0';
          WHEN "10010010110" =>
            state <= "10010010111";
            uut_rst <= '0';
          WHEN "10010010111" =>
            state <= "10010011000";
            uut_rst <= '0';
          WHEN "10010011000" =>
            state <= "10010011001";
            uut_rst <= '0';
          WHEN "10010011001" =>
            state <= "10010011010";
            uut_rst <= '0';
          WHEN "10010011010" =>
            state <= "10010011011";
            uut_rst <= '0';
          WHEN "10010011011" =>
            state <= "10010011100";
            uut_rst <= '0';
          WHEN "10010011100" =>
            state <= "10010011101";
            uut_rst <= '0';
          WHEN "10010011101" =>
            state <= "10010011110";
            uut_rst <= '0';
          WHEN "10010011110" =>
            state <= "10010011111";
            uut_rst <= '0';
          WHEN "10010011111" =>
            state <= "10010100000";
            uut_rst <= '0';
          WHEN "10010100000" =>
            state <= "10010100001";
            uut_rst <= '0';
          WHEN "10010100001" =>
            state <= "10010100010";
            uut_rst <= '0';
          WHEN "10010100010" =>
            state <= "10010100011";
            uut_rst <= '0';
          WHEN "10010100011" =>
            state <= "10010100100";
            uut_rst <= '0';
          WHEN "10010100100" =>
            state <= "10010100101";
            uut_rst <= '0';
          WHEN "10010100101" =>
            state <= "10010100110";
            uut_rst <= '0';
          WHEN "10010100110" =>
            state <= "10010100111";
            uut_rst <= '0';
          WHEN "10010100111" =>
            state <= "10010101000";
            uut_rst <= '0';
          WHEN "10010101000" =>
            state <= "10010101001";
            uut_rst <= '0';
          WHEN "10010101001" =>
            state <= "10010101010";
            uut_rst <= '0';
          WHEN "10010101010" =>
            state <= "10010101011";
            uut_rst <= '0';
          WHEN "10010101011" =>
            state <= "10010101100";
            uut_rst <= '0';
          WHEN "10010101100" =>
            state <= "10010101101";
            uut_rst <= '0';
          WHEN "10010101101" =>
            state <= "10010101110";
            uut_rst <= '0';
          WHEN "10010101110" =>
            state <= "10010101111";
            uut_rst <= '0';
          WHEN "10010101111" =>
            state <= "10010110000";
            uut_rst <= '0';
          WHEN "10010110000" =>
            state <= "10010110001";
            uut_rst <= '0';
          WHEN "10010110001" =>
            state <= "10010110010";
            uut_rst <= '0';
          WHEN "10010110010" =>
            state <= "10010110011";
            uut_rst <= '0';
          WHEN "10010110011" =>
            state <= "10010110100";
            uut_rst <= '0';
          WHEN "10010110100" =>
            state <= "10010110101";
            uut_rst <= '0';
          WHEN "10010110101" =>
            state <= "10010110110";
            uut_rst <= '0';
          WHEN "10010110110" =>
            state <= "10010110111";
            uut_rst <= '0';
          WHEN "10010110111" =>
            state <= "10010111000";
            uut_rst <= '0';
          WHEN "10010111000" =>
            state <= "10010111001";
            uut_rst <= '0';
          WHEN "10010111001" =>
            state <= "10010111010";
            uut_rst <= '0';
          WHEN "10010111010" =>
            state <= "10010111011";
            uut_rst <= '0';
          WHEN "10010111011" =>
            state <= "10010111100";
            uut_rst <= '0';
          WHEN "10010111100" =>
            state <= "10010111101";
            uut_rst <= '0';
          WHEN "10010111101" =>
            state <= "10010111110";
            uut_rst <= '0';
          WHEN "10010111110" =>
            state <= "10010111111";
            uut_rst <= '0';
          WHEN "10010111111" =>
            state <= "10011000000";
            uut_rst <= '0';
          WHEN "10011000000" =>
            state <= "10011000001";
            uut_rst <= '0';
          WHEN "10011000001" =>
            state <= "10011000010";
            uut_rst <= '0';
          WHEN "10011000010" =>
            state <= "10011000011";
            uut_rst <= '0';
          WHEN "10011000011" =>
            state <= "10011000100";
            uut_rst <= '0';
          WHEN "10011000100" =>
            state <= "10011000101";
            uut_rst <= '0';
          WHEN "10011000101" =>
            state <= "10011000110";
            uut_rst <= '0';
          WHEN "10011000110" =>
            state <= "10011000111";
            uut_rst <= '0';
          WHEN "10011000111" =>
            state <= "10011001000";
            uut_rst <= '0';
          WHEN "10011001000" =>
            state <= "10011001001";
            uut_rst <= '0';
          WHEN "10011001001" =>
            state <= "10011001010";
            uut_rst <= '0';
          WHEN "10011001010" =>
            state <= "10011001011";
            uut_rst <= '0';
          WHEN "10011001011" =>
            state <= "10011001100";
            uut_rst <= '0';
          WHEN "10011001100" =>
            state <= "10011001101";
            uut_rst <= '0';
          WHEN "10011001101" =>
            state <= "10011001110";
            uut_rst <= '0';
          WHEN "10011001110" =>
            state <= "10011001111";
            uut_rst <= '0';
          WHEN "10011001111" =>
            state <= "10011010000";
            uut_rst <= '0';
          WHEN "10011010000" =>
            state <= "10011010001";
            uut_rst <= '0';
          WHEN "10011010001" =>
            state <= "10011010010";
            uut_rst <= '0';
          WHEN "10011010010" =>
            state <= "10011010011";
            uut_rst <= '0';
          WHEN "10011010011" =>
            state <= "10011010100";
            uut_rst <= '0';
          WHEN "10011010100" =>
            state <= "10011010101";
            uut_rst <= '0';
          WHEN "10011010101" =>
            state <= "10011010110";
            uut_rst <= '0';
          WHEN "10011010110" =>
            state <= "10011010111";
            uut_rst <= '0';
          WHEN "10011010111" =>
            state <= "10011011000";
            uut_rst <= '0';
          WHEN "10011011000" =>
            state <= "10011011001";
            uut_rst <= '0';
          WHEN "10011011001" =>
            state <= "10011011010";
            uut_rst <= '0';
          WHEN "10011011010" =>
            state <= "10011011011";
            uut_rst <= '0';
          WHEN "10011011011" =>
            state <= "10011011100";
            uut_rst <= '0';
          WHEN "10011011100" =>
            state <= "10011011101";
            uut_rst <= '0';
          WHEN "10011011101" =>
            state <= "10011011110";
            uut_rst <= '0';
          WHEN "10011011110" =>
            state <= "10011011111";
            uut_rst <= '0';
          WHEN "10011011111" =>
            state <= "10011100000";
            uut_rst <= '0';
          WHEN "10011100000" =>
            state <= "10011100001";
            uut_rst <= '0';
          WHEN "10011100001" =>
            state <= "10011100010";
            uut_rst <= '0';
          WHEN "10011100010" =>
            state <= "10011100011";
            uut_rst <= '0';
          WHEN "10011100011" =>
            state <= "10011100100";
            uut_rst <= '0';
          WHEN "10011100100" =>
            state <= "10011100101";
            uut_rst <= '0';
          WHEN "10011100101" =>
            state <= "10011100110";
            uut_rst <= '0';
          WHEN "10011100110" =>
            state <= "10011100111";
            uut_rst <= '0';
          WHEN "10011100111" =>
            state <= "10011101000";
            uut_rst <= '0';
          WHEN "10011101000" =>
            state <= "10011101001";
            uut_rst <= '0';
          WHEN "10011101001" =>
            state <= "10011101010";
            uut_rst <= '0';
          WHEN "10011101010" =>
            state <= "10011101011";
            uut_rst <= '0';
          WHEN "10011101011" =>
            state <= "10011101100";
            uut_rst <= '0';
          WHEN "10011101100" =>
            state <= "10011101101";
            uut_rst <= '0';
          WHEN "10011101101" =>
            state <= "10011101110";
            uut_rst <= '0';
          WHEN "10011101110" =>
            state <= "10011101111";
            uut_rst <= '0';
          WHEN "10011101111" =>
            state <= "10011110000";
            uut_rst <= '0';
          WHEN "10011110000" =>
            state <= "10011110001";
            uut_rst <= '0';
          WHEN "10011110001" =>
            state <= "10011110010";
            uut_rst <= '0';
          WHEN "10011110010" =>
            state <= "10011110011";
            uut_rst <= '0';
          WHEN "10011110011" =>
            state <= "10011110100";
            uut_rst <= '0';
          WHEN "10011110100" =>
            state <= "10011110101";
            uut_rst <= '0';
          WHEN "10011110101" =>
            state <= "10011110110";
            uut_rst <= '0';
          WHEN "10011110110" =>
            state <= "10011110111";
            uut_rst <= '0';
          WHEN "10011110111" =>
            state <= "10011111000";
            uut_rst <= '0';
          WHEN "10011111000" =>
            state <= "10011111001";
            uut_rst <= '0';
          WHEN "10011111001" =>
            state <= "10011111010";
            uut_rst <= '0';
          WHEN "10011111010" =>
            state <= "10011111011";
            uut_rst <= '0';
          WHEN "10011111011" =>
            state <= "10011111100";
            uut_rst <= '0';
          WHEN "10011111100" =>
            state <= "10011111101";
            uut_rst <= '0';
          WHEN "10011111101" =>
            state <= "10011111110";
            uut_rst <= '0';
          WHEN "10011111110" =>
            state <= "10011111111";
            uut_rst <= '0';
          WHEN "10011111111" =>
            state <= "10100000000";
            uut_rst <= '0';
          WHEN "10100000000" =>
            state <= "10100000001";
            uut_rst <= '0';
          WHEN "10100000001" =>
            state <= "10100000010";
            uut_rst <= '0';
          WHEN "10100000010" =>
            state <= "10100000011";
            uut_rst <= '0';
          WHEN "10100000011" =>
            state <= "10100000100";
            uut_rst <= '0';
          WHEN "10100000100" =>
            state <= "10100000101";
            uut_rst <= '0';
          WHEN "10100000101" =>
            state <= "10100000110";
            uut_rst <= '0';
          WHEN "10100000110" =>
            state <= "10100000111";
            uut_rst <= '0';
          WHEN "10100000111" =>
            state <= "10100001000";
            uut_rst <= '0';
          WHEN "10100001000" =>
            state <= "10100001001";
            uut_rst <= '0';
          WHEN "10100001001" =>
            state <= "10100001010";
            uut_rst <= '0';
          WHEN "10100001010" =>
            state <= "10100001011";
            uut_rst <= '0';
          WHEN "10100001011" =>
            state <= "10100001100";
            uut_rst <= '0';
          WHEN "10100001100" =>
            state <= "10100001101";
            uut_rst <= '0';
          WHEN "10100001101" =>
            state <= "10100001110";
            uut_rst <= '0';
          WHEN "10100001110" =>
            state <= "10100001111";
            uut_rst <= '0';
          WHEN "10100001111" =>
            state <= "10100010000";
            uut_rst <= '0';
          WHEN "10100010000" =>
            state <= "10100010001";
            uut_rst <= '0';
          WHEN "10100010001" =>
            state <= "10100010010";
            uut_rst <= '0';
          WHEN "10100010010" =>
            state <= "10100010011";
            uut_rst <= '0';
          WHEN "10100010011" =>
            state <= "10100010100";
            uut_rst <= '0';
          WHEN "10100010100" =>
            state <= "10100010101";
            uut_rst <= '0';
          WHEN "10100010101" =>
            state <= "10100010110";
            uut_rst <= '0';
          WHEN "10100010110" =>
            state <= "10100010111";
            uut_rst <= '0';
          WHEN "10100010111" =>
            state <= "10100011000";
            uut_rst <= '0';
          WHEN "10100011000" =>
            state <= "10100011001";
            uut_rst <= '0';
          WHEN "10100011001" =>
            state <= "10100011010";
            uut_rst <= '0';
          WHEN "10100011010" =>
            state <= "10100011011";
            uut_rst <= '0';
          WHEN "10100011011" =>
            state <= "10100011100";
            uut_rst <= '0';
          WHEN "10100011100" =>
            state <= "10100011101";
            uut_rst <= '0';
          WHEN "10100011101" =>
            state <= "10100011110";
            uut_rst <= '0';
          WHEN "10100011110" =>
            state <= "10100011111";
            uut_rst <= '0';
          WHEN "10100011111" =>
            state <= "10100100000";
            uut_rst <= '0';
          WHEN "10100100000" =>
            state <= "10100100001";
            uut_rst <= '0';
          WHEN "10100100001" =>
            state <= "10100100010";
            uut_rst <= '0';
          WHEN "10100100010" =>
            state <= "10100100011";
            uut_rst <= '0';
          WHEN "10100100011" =>
            state <= "10100100100";
            uut_rst <= '0';
          WHEN "10100100100" =>
            state <= "10100100101";
            uut_rst <= '0';
          WHEN "10100100101" =>
            state <= "10100100110";
            uut_rst <= '0';
          WHEN "10100100110" =>
            state <= "10100100111";
            uut_rst <= '0';
          WHEN "10100100111" =>
            state <= "10100101000";
            uut_rst <= '0';
          WHEN "10100101000" =>
            state <= "10100101001";
            uut_rst <= '0';
          WHEN "10100101001" =>
            state <= "10100101010";
            uut_rst <= '0';
          WHEN "10100101010" =>
            state <= "10100101011";
            uut_rst <= '0';
          WHEN "10100101011" =>
            state <= "10100101100";
            uut_rst <= '0';
          WHEN "10100101100" =>
            state <= "10100101101";
            uut_rst <= '0';
          WHEN "10100101101" =>
            state <= "10100101110";
            uut_rst <= '0';
          WHEN "10100101110" =>
            state <= "10100101111";
            uut_rst <= '0';
          WHEN "10100101111" =>
            state <= "10100110000";
            uut_rst <= '0';
          WHEN "10100110000" =>
            state <= "10100110001";
            uut_rst <= '0';
          WHEN "10100110001" =>
            state <= "10100110010";
            uut_rst <= '0';
          WHEN "10100110010" =>
            state <= "10100110011";
            uut_rst <= '0';
          WHEN "10100110011" =>
            state <= "10100110100";
            uut_rst <= '0';
          WHEN "10100110100" =>
            state <= "10100110101";
            uut_rst <= '0';
          WHEN "10100110101" =>
            state <= "10100110110";
            uut_rst <= '0';
          WHEN "10100110110" =>
            state <= "10100110111";
            uut_rst <= '0';
          WHEN "10100110111" =>
            state <= "10100111000";
            uut_rst <= '0';
          WHEN "10100111000" =>
            state <= "10100111001";
            uut_rst <= '0';
          WHEN "10100111001" =>
            state <= "10100111010";
            uut_rst <= '0';
          WHEN "10100111010" =>
            state <= "10100111011";
            uut_rst <= '0';
          WHEN "10100111011" =>
            state <= "10100111100";
            uut_rst <= '0';
          WHEN "10100111100" =>
            state <= "10100111101";
            uut_rst <= '0';
          WHEN "10100111101" =>
            state <= "10100111110";
            uut_rst <= '0';
          WHEN "10100111110" =>
            state <= "10100111111";
            uut_rst <= '0';
          WHEN "10100111111" =>
            state <= "10101000000";
            uut_rst <= '0';
          WHEN "10101000000" =>
            state <= "10101000001";
            uut_rst <= '0';
          WHEN "10101000001" =>
            state <= "10101000010";
            uut_rst <= '0';
          WHEN "10101000010" =>
            state <= "10101000011";
            uut_rst <= '0';
          WHEN "10101000011" =>
            state <= "10101000100";
            uut_rst <= '0';
          WHEN "10101000100" =>
            state <= "10101000101";
            uut_rst <= '0';
          WHEN "10101000101" =>
            state <= "10101000110";
            uut_rst <= '0';
          WHEN "10101000110" =>
            state <= "10101000111";
            uut_rst <= '0';
          WHEN "10101000111" =>
            state <= "10101001000";
            uut_rst <= '0';
          WHEN "10101001000" =>
            state <= "10101001001";
            uut_rst <= '0';
          WHEN "10101001001" =>
            state <= "10101001010";
            uut_rst <= '0';
          WHEN "10101001010" =>
            state <= "10101001011";
            uut_rst <= '0';
          WHEN "10101001011" =>
            state <= "10101001100";
            uut_rst <= '0';
          WHEN "10101001100" =>
            state <= "10101001101";
            uut_rst <= '0';
          WHEN "10101001101" =>
            state <= "10101001110";
            uut_rst <= '0';
          WHEN "10101001110" =>
            state <= "10101001111";
            uut_rst <= '0';
          WHEN "10101001111" =>
            state <= "10101010000";
            uut_rst <= '0';
          WHEN "10101010000" =>
            state <= "10101010001";
            uut_rst <= '0';
          WHEN "10101010001" =>
            state <= "10101010010";
            uut_rst <= '0';
          WHEN "10101010010" =>
            state <= "10101010011";
            uut_rst <= '0';
          WHEN "10101010011" =>
            state <= "10101010100";
            uut_rst <= '0';
          WHEN "10101010100" =>
            state <= "10101010101";
            uut_rst <= '0';
          WHEN "10101010101" =>
            state <= "10101010110";
            uut_rst <= '0';
          WHEN "10101010110" =>
            state <= "10101010111";
            uut_rst <= '0';
          WHEN "10101010111" =>
            state <= "10101011000";
            uut_rst <= '0';
          WHEN "10101011000" =>
            state <= "10101011001";
            uut_rst <= '0';
          WHEN "10101011001" =>
            state <= "10101011010";
            uut_rst <= '0';
          WHEN "10101011010" =>
            state <= "10101011011";
            uut_rst <= '0';
          WHEN "10101011011" =>
            state <= "10101011100";
            uut_rst <= '0';
          WHEN "10101011100" =>
            state <= "10101011101";
            uut_rst <= '0';
          WHEN "10101011101" =>
            state <= "10101011110";
            uut_rst <= '0';
          WHEN "10101011110" =>
            state <= "10101011111";
            uut_rst <= '0';
          WHEN "10101011111" =>
            state <= "10101100000";
            uut_rst <= '0';
          WHEN "10101100000" =>
            state <= "10101100001";
            uut_rst <= '0';
          WHEN "10101100001" =>
            state <= "10101100010";
            uut_rst <= '0';
          WHEN "10101100010" =>
            state <= "10101100011";
            uut_rst <= '0';
          WHEN "10101100011" =>
            state <= "10101100100";
            uut_rst <= '0';
          WHEN "10101100100" =>
            state <= "10101100101";
            uut_rst <= '0';
          WHEN "10101100101" =>
            state <= "10101100110";
            uut_rst <= '0';
          WHEN "10101100110" =>
            state <= "10101100111";
            uut_rst <= '0';
          WHEN "10101100111" =>
            state <= "10101101000";
            uut_rst <= '0';
          WHEN "10101101000" =>
            state <= "10101101001";
            uut_rst <= '0';
          WHEN "10101101001" =>
            state <= "10101101010";
            uut_rst <= '0';
          WHEN "10101101010" =>
            state <= "10101101011";
            uut_rst <= '0';
          WHEN "10101101011" =>
            state <= "10101101100";
            uut_rst <= '0';
          WHEN "10101101100" =>
            state <= "10101101101";
            uut_rst <= '0';
          WHEN "10101101101" =>
            state <= "10101101110";
            uut_rst <= '0';
          WHEN "10101101110" =>
            state <= "10101101111";
            uut_rst <= '0';
          WHEN "10101101111" =>
            state <= "10101110000";
            uut_rst <= '0';
          WHEN "10101110000" =>
            state <= "10101110001";
            uut_rst <= '0';
          WHEN "10101110001" =>
            state <= "10101110010";
            uut_rst <= '0';
          WHEN "10101110010" =>
            state <= "10101110011";
            uut_rst <= '0';
          WHEN "10101110011" =>
            state <= "10101110100";
            uut_rst <= '0';
          WHEN "10101110100" =>
            state <= "10101110101";
            uut_rst <= '0';
          WHEN "10101110101" =>
            state <= "10101110110";
            uut_rst <= '0';
          WHEN "10101110110" =>
            state <= "10101110111";
            uut_rst <= '0';
          WHEN "10101110111" =>
            state <= "10101111000";
            uut_rst <= '0';
          WHEN "10101111000" =>
            state <= "10101111001";
            uut_rst <= '0';
          WHEN "10101111001" =>
            state <= "10101111010";
            uut_rst <= '0';
          WHEN "10101111010" =>
            state <= "10101111011";
            uut_rst <= '0';
          WHEN "10101111011" =>
            state <= "10101111100";
            uut_rst <= '0';
          WHEN "10101111100" =>
            state <= "10101111101";
            uut_rst <= '0';
          WHEN "10101111101" =>
            state <= "10101111110";
            uut_rst <= '0';
          WHEN "10101111110" =>
            state <= "10101111111";
            uut_rst <= '0';
          WHEN "10101111111" =>
            state <= "10110000000";
            uut_rst <= '0';
          WHEN "10110000000" =>
            state <= "10110000001";
            uut_rst <= '0';
          WHEN "10110000001" =>
            state <= "10110000010";
            uut_rst <= '0';
          WHEN "10110000010" =>
            state <= "10110000011";
            uut_rst <= '0';
          WHEN "10110000011" =>
            state <= "10110000100";
            uut_rst <= '0';
          WHEN "10110000100" =>
            state <= "10110000101";
            uut_rst <= '0';
          WHEN "10110000101" =>
            state <= "10110000110";
            uut_rst <= '0';
          WHEN "10110000110" =>
            state <= "10110000111";
            uut_rst <= '0';
          WHEN "10110000111" =>
            state <= "10110001000";
            uut_rst <= '0';
          WHEN "10110001000" =>
            state <= "10110001001";
            uut_rst <= '0';
          WHEN "10110001001" =>
            state <= "10110001010";
            uut_rst <= '0';
          WHEN "10110001010" =>
            state <= "10110001011";
            uut_rst <= '0';
          WHEN "10110001011" =>
            state <= "10110001100";
            uut_rst <= '0';
          WHEN "10110001100" =>
            state <= "10110001101";
            uut_rst <= '0';
          WHEN "10110001101" =>
            state <= "10110001110";
            uut_rst <= '0';
          WHEN "10110001110" =>
            state <= "10110001111";
            uut_rst <= '0';
          WHEN "10110001111" =>
            state <= "10110010000";
            uut_rst <= '0';
          WHEN "10110010000" =>
            state <= "10110010001";
            uut_rst <= '0';
          WHEN "10110010001" =>
            state <= "10110010010";
            uut_rst <= '0';
          WHEN "10110010010" =>
            state <= "10110010011";
            uut_rst <= '0';
          WHEN "10110010011" =>
            state <= "10110010100";
            uut_rst <= '0';
          WHEN "10110010100" =>
            state <= "10110010101";
            uut_rst <= '0';
          WHEN "10110010101" =>
            state <= "10110010110";
            uut_rst <= '0';
          WHEN "10110010110" =>
            state <= "10110010111";
            uut_rst <= '0';
          WHEN "10110010111" =>
            state <= "10110011000";
            uut_rst <= '0';
          WHEN "10110011000" =>
            state <= "10110011001";
            uut_rst <= '0';
          WHEN "10110011001" =>
            state <= "10110011010";
            uut_rst <= '0';
          WHEN "10110011010" =>
            state <= "10110011011";
            uut_rst <= '0';
          WHEN "10110011011" =>
            state <= "10110011100";
            uut_rst <= '0';
          WHEN "10110011100" =>
            state <= "10110011101";
            uut_rst <= '0';
          WHEN "10110011101" =>
            state <= "10110011110";
            uut_rst <= '0';
          WHEN "10110011110" =>
            state <= "10110011111";
            uut_rst <= '0';
          WHEN "10110011111" =>
            state <= "10110100000";
            uut_rst <= '0';
          WHEN "10110100000" =>
            state <= "10110100001";
            uut_rst <= '0';
          WHEN "10110100001" =>
            state <= "10110100010";
            uut_rst <= '0';
          WHEN "10110100010" =>
            state <= "10110100011";
            uut_rst <= '0';
          WHEN "10110100011" =>
            state <= "10110100100";
            uut_rst <= '0';
          WHEN "10110100100" =>
            state <= "10110100101";
            uut_rst <= '0';
          WHEN "10110100101" =>
            state <= "10110100110";
            uut_rst <= '0';
          WHEN "10110100110" =>
            state <= "10110100111";
            uut_rst <= '0';
          WHEN "10110100111" =>
            state <= "10110101000";
            uut_rst <= '0';
          WHEN "10110101000" =>
            state <= "10110101001";
            uut_rst <= '0';
          WHEN "10110101001" =>
            state <= "10110101010";
            uut_rst <= '0';
          WHEN "10110101010" =>
            state <= "10110101011";
            uut_rst <= '0';
          WHEN "10110101011" =>
            state <= "10110101100";
            uut_rst <= '0';
          WHEN "10110101100" =>
            state <= "10110101101";
            uut_rst <= '0';
          WHEN "10110101101" =>
            state <= "10110101110";
            uut_rst <= '0';
          WHEN "10110101110" =>
            state <= "10110101111";
            uut_rst <= '0';
          WHEN "10110101111" =>
            state <= "10110110000";
            uut_rst <= '0';
          WHEN "10110110000" =>
            state <= "10110110001";
            uut_rst <= '0';
          WHEN "10110110001" =>
            state <= "10110110010";
            uut_rst <= '0';
          WHEN "10110110010" =>
            state <= "10110110011";
            uut_rst <= '0';
          WHEN "10110110011" =>
            state <= "10110110100";
            uut_rst <= '0';
          WHEN "10110110100" =>
            state <= "10110110101";
            uut_rst <= '0';
          WHEN "10110110101" =>
            state <= "10110110110";
            uut_rst <= '0';
          WHEN "10110110110" =>
            state <= "10110110111";
            uut_rst <= '0';
          WHEN "10110110111" =>
            state <= "10110111000";
            uut_rst <= '0';
          WHEN "10110111000" =>
            state <= "10110111001";
            uut_rst <= '0';
          WHEN "10110111001" =>
            state <= "10110111010";
            uut_rst <= '0';
          WHEN "10110111010" =>
            state <= "10110111011";
            uut_rst <= '0';
          WHEN "10110111011" =>
            state <= "10110111100";
            uut_rst <= '0';
          WHEN "10110111100" =>
            state <= "10110111101";
            uut_rst <= '0';
          WHEN "10110111101" =>
            state <= "10110111110";
            uut_rst <= '0';
          WHEN "10110111110" =>
            state <= "10110111111";
            uut_rst <= '0';
          WHEN "10110111111" =>
            state <= "10111000000";
            uut_rst <= '0';
          WHEN "10111000000" =>
            state <= "10111000001";
            uut_rst <= '0';
          WHEN "10111000001" =>
            state <= "10111000010";
            uut_rst <= '0';
          WHEN "10111000010" =>
            state <= "10111000011";
            uut_rst <= '0';
          WHEN "10111000011" =>
            state <= "10111000100";
            uut_rst <= '0';
          WHEN "10111000100" =>
            state <= "10111000101";
            uut_rst <= '0';
          WHEN "10111000101" =>
            state <= "10111000110";
            uut_rst <= '0';
          WHEN "10111000110" =>
            state <= "10111000111";
            uut_rst <= '0';
          WHEN "10111000111" =>
            state <= "10111001000";
            uut_rst <= '0';
          WHEN "10111001000" =>
            state <= "10111001001";
            uut_rst <= '0';
          WHEN "10111001001" =>
            state <= "10111001010";
            uut_rst <= '0';
          WHEN "10111001010" =>
            state <= "10111001011";
            uut_rst <= '0';
          WHEN "10111001011" =>
            state <= "10111001100";
            uut_rst <= '0';
          WHEN "10111001100" =>
            state <= "10111001101";
            uut_rst <= '0';
          WHEN "10111001101" =>
            state <= "10111001110";
            uut_rst <= '0';
          WHEN "10111001110" =>
            state <= "10111001111";
            uut_rst <= '0';
          WHEN "10111001111" =>
            state <= "10111010000";
            uut_rst <= '0';
          WHEN "10111010000" =>
            state <= "10111010001";
            uut_rst <= '0';
          WHEN "10111010001" =>
            state <= "10111010010";
            uut_rst <= '0';
          WHEN "10111010010" =>
            state <= "10111010011";
            uut_rst <= '0';
          WHEN "10111010011" =>
            state <= "10111010100";
            uut_rst <= '0';
          WHEN "10111010100" =>
            state <= "10111010101";
            uut_rst <= '0';
          WHEN "10111010101" =>
            state <= "10111010110";
            uut_rst <= '0';
          WHEN "10111010110" =>
            state <= "10111010111";
            uut_rst <= '0';
          WHEN "10111010111" =>
            state <= "10111011000";
            uut_rst <= '0';
          WHEN "10111011000" =>
            state <= "10111011001";
            uut_rst <= '0';
          WHEN "10111011001" =>
            state <= "10111011010";
            uut_rst <= '0';
          WHEN "10111011010" =>
            state <= "10111011011";
            uut_rst <= '0';
          WHEN "10111011011" =>
            state <= "10111011100";
            uut_rst <= '0';
          WHEN "10111011100" =>
            state <= "10111011101";
            uut_rst <= '0';
          WHEN "10111011101" =>
            state <= "10111011110";
            uut_rst <= '0';
          WHEN "10111011110" =>
            state <= "10111011111";
            uut_rst <= '0';
          WHEN "10111011111" =>
            state <= "10111100000";
            uut_rst <= '0';
          WHEN "10111100000" =>
            state <= "10111100001";
            uut_rst <= '0';
          WHEN "10111100001" =>
            state <= "10111100010";
            uut_rst <= '0';
          WHEN "10111100010" =>
            state <= "10111100011";
            uut_rst <= '0';
          WHEN "10111100011" =>
            state <= "10111100100";
            uut_rst <= '0';
          WHEN "10111100100" =>
            state <= "10111100101";
            uut_rst <= '0';
          WHEN "10111100101" =>
            state <= "10111100110";
            uut_rst <= '0';
          WHEN "10111100110" =>
            state <= "10111100111";
            uut_rst <= '0';
          WHEN "10111100111" =>
            state <= "10111101000";
            uut_rst <= '0';
          WHEN "10111101000" =>
            state <= "10111101001";
            uut_rst <= '0';
          WHEN "10111101001" =>
            state <= "10111101010";
            uut_rst <= '0';
          WHEN "10111101010" =>
            state <= "10111101011";
            uut_rst <= '0';
          WHEN "10111101011" =>
            state <= "10111101100";
            uut_rst <= '0';
          WHEN "10111101100" =>
            state <= "10111101101";
            uut_rst <= '0';
          WHEN "10111101101" =>
            state <= "10111101110";
            uut_rst <= '0';
          WHEN "10111101110" =>
            state <= "10111101111";
            uut_rst <= '0';
          WHEN "10111101111" =>
            state <= "10111110000";
            uut_rst <= '0';
          WHEN "10111110000" =>
            state <= "10111110001";
            uut_rst <= '0';
          WHEN "10111110001" =>
            state <= "10111110010";
            uut_rst <= '0';
          WHEN "10111110010" =>
            state <= "10111110011";
            uut_rst <= '0';
          WHEN "10111110011" =>
            state <= "10111110100";
            uut_rst <= '0';
          WHEN "10111110100" =>
            state <= "10111110101";
            uut_rst <= '0';
          WHEN "10111110101" =>
            state <= "10111110110";
            uut_rst <= '0';
          WHEN "10111110110" =>
            state <= "10111110111";
            uut_rst <= '0';
          WHEN "10111110111" =>
            state <= "10111111000";
            uut_rst <= '0';
          WHEN "10111111000" =>
            state <= "10111111001";
            uut_rst <= '0';
          WHEN "10111111001" =>
            state <= "10111111010";
            uut_rst <= '0';
          WHEN "10111111010" =>
            state <= "10111111011";
            uut_rst <= '0';
          WHEN "10111111011" =>
            state <= "10111111100";
            uut_rst <= '0';
          WHEN "10111111100" =>
            state <= "10111111101";
            uut_rst <= '0';
          WHEN "10111111101" =>
            state <= "10111111110";
            uut_rst <= '0';
          WHEN "10111111110" =>
            state <= "10111111111";
            uut_rst <= '0';
          WHEN "10111111111" =>
            state <= "11000000000";
            uut_rst <= '0';
          WHEN "11000000000" =>
            state <= "11000000001";
            uut_rst <= '0';
          WHEN "11000000001" =>
            state <= "11000000010";
            uut_rst <= '0';
          WHEN "11000000010" =>
            state <= "11000000011";
            uut_rst <= '0';
          WHEN "11000000011" =>
            state <= "11000000100";
            uut_rst <= '0';
          WHEN "11000000100" =>
            state <= "11000000101";
            uut_rst <= '0';
          WHEN "11000000101" =>
            state <= "11000000110";
            uut_rst <= '0';
          WHEN "11000000110" =>
            state <= "11000000111";
            uut_rst <= '0';
          WHEN "11000000111" =>
            state <= "11000001000";
            uut_rst <= '0';
          WHEN "11000001000" =>
            state <= "11000001001";
            uut_rst <= '0';
          WHEN "11000001001" =>
            state <= "11000001010";
            uut_rst <= '0';
          WHEN "11000001010" =>
            state <= "11000001011";
            uut_rst <= '0';
          WHEN "11000001011" =>
            state <= "11000001100";
            uut_rst <= '0';
          WHEN "11000001100" =>
            state <= "11000001101";
            uut_rst <= '0';
          WHEN "11000001101" =>
            state <= "11000001110";
            uut_rst <= '0';
          WHEN "11000001110" =>
            state <= "11000001111";
            uut_rst <= '0';
          WHEN "11000001111" =>
            state <= "11000010000";
            uut_rst <= '0';
          WHEN "11000010000" =>
            state <= "11000010001";
            uut_rst <= '0';
          WHEN "11000010001" =>
            state <= "11000010010";
            uut_rst <= '0';
          WHEN "11000010010" =>
            state <= "11000010011";
            uut_rst <= '0';
          WHEN OTHERS =>
            DONE <= '1';
            uut_rst <= '1';
        END CASE;
      END IF;
    END IF;
  END PROCESS;
END;
