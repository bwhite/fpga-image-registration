-- Module Name:  i2c_core.vhd
-- File Description:  Generic i2c module with write capability only.
-- Project:  FPGA Image Registration
-- Target Device:  XC5VSX50T (Xilinx Virtex5 SXT)
-- Target Board:  ML506
-- Synthesis Tool:  Xilinx ISE 9.2
-- Copyright (C) 2008 Brandyn Allen White
-- Contact:  bwhite(at)cs.ucf.edu
-- Project Website:  http://code.google.com/p/fpga-image-registration/

-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.

-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the
-- GNU General Public License for more details.

-- You should have received a copy of the GNU General Public License
-- along with this program. If not, see <http://www.gnu.org/licenses/>.

-- NOTE The data is in little endian byte ordering, data is sent lowest byte
-- first, highest bit first (I2C convention).

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


ENTITY i2c_core IS
  PORT (clk           : IN  std_logic;
        data          : IN  std_logic_vector (23 DOWNTO 0);
        new_data      : IN  std_logic;
        reset         : IN  std_logic;
        i2c_sda       : OUT std_logic;
        i2c_scl       : OUT std_logic;
        received_data : OUT std_logic);
END i2c_core;

ARCHITECTURE Behavioral OF i2c_core IS
  SIGNAL cur_data          : std_logic_vector (23 DOWNTO 0);  -- {device_id(7 downto 0), address(7 downto 0), data(7 downto 0)}
  SIGNAL i2c_state         : std_logic_vector (2 DOWNTO 0) := (OTHERS => '0');  -- {START, DATA, POST_DATA, STOP, STOP_WAIT, X, X, X}
  SIGNAL byte_position     : std_logic_vector(1 DOWNTO 0)  := (OTHERS => '0');  -- {device_id, address, data, X}
  SIGNAL bit_position      : std_logic_vector(2 DOWNTO 0)  := (OTHERS => '0');
  SIGNAL received_data_reg : std_logic                     := '0';
  SIGNAL i2c_sda_reg       : std_logic                     := '1';

-- I2C Clock Variables
  SIGNAL i2c_clock_counter    : std_logic_vector (8 DOWNTO 0) := (OTHERS => '0');  -- [0,499]
  SIGNAL i2c_edge_count       : std_logic_vector (2 DOWNTO 0) := (OTHERS => '0');  -- [0,4]
  SIGNAL i2c_clock            : std_logic                     := '1';
  SIGNAL i2c_clock_5x         : std_logic                     := '1';
  SIGNAL i2c_clock_5x_posedge : std_logic                     := '1';

BEGIN
  i2c_scl       <= '0' WHEN i2c_clock = '0'   ELSE 'Z';  -- Output using {0,Z logic}
  i2c_sda       <= '0' WHEN i2c_sda_reg = '0' ELSE 'Z';  -- Output using {0,Z logic}
  received_data <= received_data_reg;

  PROCESS(clk)
  BEGIN
    IF (clk'event AND clk = '1') THEN
      -- Set initial register values upon synchronous reset
      IF (reset = '1') THEN
        i2c_state         <= (OTHERS => '0');
        byte_position     <= (OTHERS => '0');
        bit_position      <= (OTHERS => '0');
        received_data_reg <= '0';
        i2c_sda_reg       <= '1';

        -- I2C Clock Variables
        i2c_clock_counter    <= (OTHERS => '0');
        i2c_edge_count       <= (OTHERS => '0');
        i2c_clock            <= '1';
        i2c_clock_5x         <= '1';
        i2c_clock_5x_posedge <= '1';
      ELSE
        -- If we are supposed to start; however, no data is ready, then reset the clock logic to hold it high
        IF (i2c_state = "000" AND new_data = '0') THEN
          i2c_sda_reg       <= '1';
          received_data_reg <= '0';

                                        -- I2C Clock Variables
          i2c_clock_counter    <= (OTHERS => '0');
          i2c_edge_count       <= (OTHERS => '0');
          i2c_clock            <= '1';
          i2c_clock_5x         <= '1';
          i2c_clock_5x_posedge <= '1';
        ELSE
                                        -- I2C Clock generation - Reduces clock rate by 100 for internal use and 500 for external use.
          IF (i2c_clock_counter = 99 OR i2c_clock_counter = 199 OR i2c_clock_counter = 299 OR i2c_clock_counter = 399 OR i2c_clock_counter = 499) THEN
            i2c_clock_5x <= NOT i2c_clock_5x;
            IF (i2c_clock_5x = '0') THEN
              i2c_clock_5x_posedge <= '1';
              IF (i2c_edge_count < 4) THEN
                i2c_edge_count <= i2c_edge_count + 1;
              ELSE
                i2c_edge_count <= (OTHERS => '0');
              END IF;
            END IF;
          END IF;

                                        -- Toggle the external I2C clock every 500 ticks
          IF (i2c_clock_counter = 499) THEN
            i2c_clock_counter <= (OTHERS => '0');
            i2c_clock         <= NOT i2c_clock;
          ELSE
            i2c_clock_counter <= i2c_clock_counter + 1;
          END IF;
        END IF;

        -- Main I2C Logic
        IF (i2c_clock_5x_posedge = '1') THEN
          i2c_clock_5x_posedge <= '0';
          CASE i2c_edge_count IS  -- Edge selection -> individual state selection
            WHEN "001" =>
              IF (i2c_state = "011") THEN      -- STATE: stop
                i2c_sda_reg <= '1';
                i2c_state   <= "000";   -- 'start'
              END IF;
            WHEN "010" =>
              IF (i2c_state = "000") THEN      -- STATE: start
                IF (new_data = '1' AND received_data_reg = '0') THEN
                  i2c_sda_reg       <= '0';
                  cur_data          <= data;
                  received_data_reg <= '1';
                  i2c_state         <= "001";  -- 'data'
                END IF;
              END IF;

            WHEN "100" =>
              CASE i2c_state IS
                WHEN "001" =>           -- STATE: data
                  CASE bit_position IS  -- Select bit position and output it (NOTE:  MSB is output first!), TODO investigate other bit selection methods
                    WHEN "000" =>
                      i2c_sda_reg <= cur_data(7);
                    WHEN "001" =>
                      i2c_sda_reg <= cur_data(6);
                    WHEN "010" =>
                      i2c_sda_reg <= cur_data(5);
                    WHEN "011" =>
                      i2c_sda_reg <= cur_data(4);
                    WHEN "100" =>
                      i2c_sda_reg <= cur_data(3);
                    WHEN "101" =>
                      i2c_sda_reg <= cur_data(2);
                    WHEN "110" =>
                      i2c_sda_reg <= cur_data(1);
                    WHEN "111" =>
                      i2c_sda_reg <= cur_data(0);
                    WHEN OTHERS =>
                      NULL;
                  END CASE;
                      bit_position <= bit_position + 1;
                      IF (bit_position = "111") THEN
                        i2c_state <= "010";  -- 'post_data'
                      ELSE
                        i2c_state <= "001";  -- 'data'
                      END IF;
                WHEN "010" =>           -- STATE: post_data
                  cur_data(15 DOWNTO 0) <= cur_data(23 DOWNTO 8);  -- Shift right by 8, TODO investigate other shifting methods
                  i2c_sda_reg           <= '1';
                  IF (byte_position = 2) THEN
                    byte_position <= (OTHERS => '0');
                    i2c_state     <= "100";
                  ELSE
                    byte_position <= byte_position + 1;
                    i2c_state     <= "001";
                  END IF;
                WHEN "100" =>           -- STATE: stop_wait
                  i2c_sda_reg <= '0';
                  i2c_state   <= "011";      -- 'stop'
                WHEN OTHERS =>
                  NULL;
              END CASE;
            WHEN OTHERS =>
              NULL;
          END CASE;
        END IF;

        -- Data synchronization acknowledgement
        IF (new_data = '0' AND received_data_reg = '1') THEN
          received_data_reg <= '0';
        END IF;
      END IF;
    END IF;
  END PROCESS;
END Behavioral;

