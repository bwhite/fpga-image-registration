/home/brandyn/fpga-image-registration/modules/./gauss_elim/div1.vhd