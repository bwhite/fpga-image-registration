/home/brandyn/fpga-image-registration/modules/./gauss_elim/div1_test.vhd