LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
ENTITY gauss_elimT0_tb IS
PORT(
  CLK : IN STD_LOGIC;
  RST : IN STD_LOGIC;
  DONE : OUT STD_LOGIC;
  FAIL : OUT STD_LOGIC;
  FAIL_NUM : OUT STD_LOGIC_VECTOR(8 DOWNTO 0));
END gauss_elimT0_tb;
ARCHITECTURE behavior OF gauss_elimT0_tb IS
  COMPONENT gauss_elim
  PORT(
    CLK : IN STD_LOGIC;
    RST : IN STD_LOGIC;
    INPUT_LOAD : IN STD_LOGIC;
    A_0_0 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_0_1 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_0_2 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_0_3 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_0_4 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_0_5 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_1_0 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_1_1 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_1_2 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_1_3 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_1_4 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_1_5 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_2_0 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_2_1 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_2_2 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_2_3 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_2_4 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_2_5 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_3_0 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_3_1 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_3_2 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_3_3 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_3_4 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_3_5 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_4_0 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_4_1 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_4_2 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_4_3 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_4_4 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_4_5 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_5_0 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_5_1 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_5_2 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_5_3 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_5_4 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_5_5 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    B_0 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    B_1 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    B_2 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    B_3 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    B_4 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    B_5 : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    X_0 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    X_1 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    X_2 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    X_3 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    X_4 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    X_5 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    OUTPUT_VALID : OUT STD_LOGIC);
  END COMPONENT;
  SIGNAL uut_rst_wire, uut_rst : STD_LOGIC;
  SIGNAL state : STD_LOGIC_VECTOR(9 DOWNTO 0);
  -- UUT Input
  SIGNAL uut_input_load : STD_LOGIC;
  SIGNAL uut_a_0_0, uut_a_0_1, uut_a_0_2, uut_a_0_3, uut_a_0_4, uut_a_0_5, uut_a_1_0, uut_a_1_1, uut_a_1_2, uut_a_1_3, uut_a_1_4, uut_a_1_5, uut_a_2_0, uut_a_2_1, uut_a_2_2, uut_a_2_3, uut_a_2_4, uut_a_2_5, uut_a_3_0, uut_a_3_1, uut_a_3_2, uut_a_3_3, uut_a_3_4, uut_a_3_5, uut_a_4_0, uut_a_4_1, uut_a_4_2, uut_a_4_3, uut_a_4_4, uut_a_4_5, uut_a_5_0, uut_a_5_1, uut_a_5_2, uut_a_5_3, uut_a_5_4, uut_a_5_5, uut_b_0, uut_b_1, uut_b_2, uut_b_3, uut_b_4, uut_b_5 : STD_LOGIC_VECTOR(26 DOWNTO 0);
  -- UUT Output
  SIGNAL uut_output_valid : STD_LOGIC;
  SIGNAL uut_x_0, uut_x_1, uut_x_2, uut_x_3, uut_x_4, uut_x_5 : STD_LOGIC_VECTOR(26 DOWNTO 0);
BEGIN
  uut_rst_wire <= RST OR uut_rst;
  uut :  gauss_elim PORT MAP (
    CLK => CLK,
    RST => uut_rst_wire,
    INPUT_LOAD => uut_input_load,
    A_0_0 => uut_a_0_0,
    A_0_1 => uut_a_0_1,
    A_0_2 => uut_a_0_2,
    A_0_3 => uut_a_0_3,
    A_0_4 => uut_a_0_4,
    A_0_5 => uut_a_0_5,
    A_1_0 => uut_a_1_0,
    A_1_1 => uut_a_1_1,
    A_1_2 => uut_a_1_2,
    A_1_3 => uut_a_1_3,
    A_1_4 => uut_a_1_4,
    A_1_5 => uut_a_1_5,
    A_2_0 => uut_a_2_0,
    A_2_1 => uut_a_2_1,
    A_2_2 => uut_a_2_2,
    A_2_3 => uut_a_2_3,
    A_2_4 => uut_a_2_4,
    A_2_5 => uut_a_2_5,
    A_3_0 => uut_a_3_0,
    A_3_1 => uut_a_3_1,
    A_3_2 => uut_a_3_2,
    A_3_3 => uut_a_3_3,
    A_3_4 => uut_a_3_4,
    A_3_5 => uut_a_3_5,
    A_4_0 => uut_a_4_0,
    A_4_1 => uut_a_4_1,
    A_4_2 => uut_a_4_2,
    A_4_3 => uut_a_4_3,
    A_4_4 => uut_a_4_4,
    A_4_5 => uut_a_4_5,
    A_5_0 => uut_a_5_0,
    A_5_1 => uut_a_5_1,
    A_5_2 => uut_a_5_2,
    A_5_3 => uut_a_5_3,
    A_5_4 => uut_a_5_4,
    A_5_5 => uut_a_5_5,
    B_0 => uut_b_0,
    B_1 => uut_b_1,
    B_2 => uut_b_2,
    B_3 => uut_b_3,
    B_4 => uut_b_4,
    B_5 => uut_b_5,
    X_0 => uut_x_0,
    X_1 => uut_x_1,
    X_2 => uut_x_2,
    X_3 => uut_x_3,
    X_4 => uut_x_4,
    X_5 => uut_x_5,
    OUTPUT_VALID => uut_output_valid
  );
  PROCESS (CLK) IS
  BEGIN
    IF CLK'event AND CLK='1' THEN
      IF RST='1' THEN
        DONE <= '0';
        FAIL <= '0';
        uut_rst <= '1';
        FAIL_NUM <= (OTHERS => '0');
        state <= (OTHERS => '0');
      ELSE
        CASE state IS
          WHEN "0000000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000000001";
            uut_rst <= '0';
          WHEN "0000000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000000010";
            uut_rst <= '0';
          WHEN "0000000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000000011";
            uut_rst <= '0';
          WHEN "0000000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000000100";
            uut_rst <= '0';
          WHEN "0000000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000000101";
            uut_rst <= '0';
          WHEN "0000000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000000110";
            uut_rst <= '0';
          WHEN "0000000110" =>
            uut_input_load <= '1';
            uut_a_0_0 <= "000000000011000011010110100";
            uut_a_0_1 <= "000000001100111111000011100";
            uut_a_0_2 <= "000000111001100101001111000";
            uut_a_0_3 <= "000000000000000010001010010";
            uut_a_0_4 <= "000000000111100110101010100";
            uut_a_0_5 <= "111111111101000110011001000";
            uut_a_1_0 <= "000000000000000110011111100";
            uut_a_1_1 <= "000000100010110101001001111";
            uut_a_1_2 <= "000000000110100011000110110";
            uut_a_1_3 <= "000000000000000011110011010";
            uut_a_1_4 <= "111111111111110101011011101";
            uut_a_1_5 <= "000000000000010010011110001";
            uut_a_2_0 <= "000000000000011100110010100";
            uut_a_2_1 <= "000000000110100011000110110";
            uut_a_2_2 <= "000000010011101111110011100";
            uut_a_2_3 <= "111111111111111110100011001";
            uut_a_2_4 <= "000000000000010010011110001";
            uut_a_2_5 <= "111111111110101101111000110";
            uut_a_3_0 <= "000000000000000010001010010";
            uut_a_3_1 <= "000000000111100110101010100";
            uut_a_3_2 <= "111111111101000110011001000";
            uut_a_3_3 <= "000000000100001110101100001";
            uut_a_3_4 <= "000001101101010011010000101";
            uut_a_3_5 <= "000000011110111111111010000";
            uut_a_4_0 <= "000000000000000011110011010";
            uut_a_4_1 <= "111111111111110101011011101";
            uut_a_4_2 <= "000000000000010010011110001";
            uut_a_4_3 <= "000000000000110110101001101";
            uut_a_4_4 <= "000001000000011100000111000";
            uut_a_4_5 <= "000000000011100110111011111";
            uut_a_5_0 <= "111111111111111110100011001";
            uut_a_5_1 <= "000000000000010010011110001";
            uut_a_5_2 <= "111111111110101101111000110";
            uut_a_5_3 <= "000000000000001111011111111";
            uut_a_5_4 <= "000000000011100110111011111";
            uut_a_5_5 <= "000000010101101100011000110";
            state <= "0000000111";
            uut_rst <= '0';
          WHEN "0000000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000001000";
            uut_rst <= '0';
          WHEN "0000001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000001001";
            uut_rst <= '0';
          WHEN "0000001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000001010";
            uut_rst <= '0';
          WHEN "0000001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000001011";
            uut_rst <= '0';
          WHEN "0000001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000001100";
            uut_rst <= '0';
          WHEN "0000001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000001101";
            uut_rst <= '0';
          WHEN "0000001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000001110";
            uut_rst <= '0';
          WHEN "0000001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000001111";
            uut_rst <= '0';
          WHEN "0000001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000010000";
            uut_rst <= '0';
          WHEN "0000010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000010001";
            uut_rst <= '0';
          WHEN "0000010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000010010";
            uut_rst <= '0';
          WHEN "0000010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000010011";
            uut_rst <= '0';
          WHEN "0000010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000010100";
            uut_rst <= '0';
          WHEN "0000010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000010101";
            uut_rst <= '0';
          WHEN "0000010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000010110";
            uut_rst <= '0';
          WHEN "0000010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000010111";
            uut_rst <= '0';
          WHEN "0000010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000011000";
            uut_rst <= '0';
          WHEN "0000011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000011001";
            uut_rst <= '0';
          WHEN "0000011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000011010";
            uut_rst <= '0';
          WHEN "0000011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000011011";
            uut_rst <= '0';
          WHEN "0000011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000011100";
            uut_rst <= '0';
          WHEN "0000011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000011101";
            uut_rst <= '0';
          WHEN "0000011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000011110";
            uut_rst <= '0';
          WHEN "0000011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000011111";
            uut_rst <= '0';
          WHEN "0000011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000100000";
            uut_rst <= '0';
          WHEN "0000100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000100001";
            uut_rst <= '0';
          WHEN "0000100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000100010";
            uut_rst <= '0';
          WHEN "0000100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000100011";
            uut_rst <= '0';
          WHEN "0000100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000100100";
            uut_rst <= '0';
          WHEN "0000100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000100101";
            uut_rst <= '0';
          WHEN "0000100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000100110";
            uut_rst <= '0';
          WHEN "0000100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000100111";
            uut_rst <= '0';
          WHEN "0000100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000101000";
            uut_rst <= '0';
          WHEN "0000101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000101001";
            uut_rst <= '0';
          WHEN "0000101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000101010";
            uut_rst <= '0';
          WHEN "0000101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000101011";
            uut_rst <= '0';
          WHEN "0000101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000101100";
            uut_rst <= '0';
          WHEN "0000101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000101101";
            uut_rst <= '0';
          WHEN "0000101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000101110";
            uut_rst <= '0';
          WHEN "0000101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000101111";
            uut_rst <= '0';
          WHEN "0000101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000110000";
            uut_rst <= '0';
          WHEN "0000110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000110001";
            uut_rst <= '0';
          WHEN "0000110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000110010";
            uut_rst <= '0';
          WHEN "0000110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000110011";
            uut_rst <= '0';
          WHEN "0000110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000110100";
            uut_rst <= '0';
          WHEN "0000110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000110101";
            uut_rst <= '0';
          WHEN "0000110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000110110";
            uut_rst <= '0';
          WHEN "0000110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000110111";
            uut_rst <= '0';
          WHEN "0000110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000111000";
            uut_rst <= '0';
          WHEN "0000111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000111001";
            uut_rst <= '0';
          WHEN "0000111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000111010";
            uut_rst <= '0';
          WHEN "0000111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000111011";
            uut_rst <= '0';
          WHEN "0000111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000111100";
            uut_rst <= '0';
          WHEN "0000111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000111101";
            uut_rst <= '0';
          WHEN "0000111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000111110";
            uut_rst <= '0';
          WHEN "0000111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0000111111";
            uut_rst <= '0';
          WHEN "0000111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001000000";
            uut_rst <= '0';
          WHEN "0001000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001000001";
            uut_rst <= '0';
          WHEN "0001000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001000010";
            uut_rst <= '0';
          WHEN "0001000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001000011";
            uut_rst <= '0';
          WHEN "0001000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001000100";
            uut_rst <= '0';
          WHEN "0001000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001000101";
            uut_rst <= '0';
          WHEN "0001000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001000110";
            uut_rst <= '0';
          WHEN "0001000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001000111";
            uut_rst <= '0';
          WHEN "0001000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001001000";
            uut_rst <= '0';
          WHEN "0001001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001001001";
            uut_rst <= '0';
          WHEN "0001001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001001010";
            uut_rst <= '0';
          WHEN "0001001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001001011";
            uut_rst <= '0';
          WHEN "0001001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001001100";
            uut_rst <= '0';
          WHEN "0001001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001001101";
            uut_rst <= '0';
          WHEN "0001001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001001110";
            uut_rst <= '0';
          WHEN "0001001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001001111";
            uut_rst <= '0';
          WHEN "0001001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001010000";
            uut_rst <= '0';
          WHEN "0001010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001010001";
            uut_rst <= '0';
          WHEN "0001010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001010010";
            uut_rst <= '0';
          WHEN "0001010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001010011";
            uut_rst <= '0';
          WHEN "0001010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001010100";
            uut_rst <= '0';
          WHEN "0001010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001010101";
            uut_rst <= '0';
          WHEN "0001010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001010110";
            uut_rst <= '0';
          WHEN "0001010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001010111";
            uut_rst <= '0';
          WHEN "0001010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001011000";
            uut_rst <= '0';
          WHEN "0001011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001011001";
            uut_rst <= '0';
          WHEN "0001011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001011010";
            uut_rst <= '0';
          WHEN "0001011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001011011";
            uut_rst <= '0';
          WHEN "0001011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001011100";
            uut_rst <= '0';
          WHEN "0001011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001011101";
            uut_rst <= '0';
          WHEN "0001011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001011110";
            uut_rst <= '0';
          WHEN "0001011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001011111";
            uut_rst <= '0';
          WHEN "0001011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001100000";
            uut_rst <= '0';
          WHEN "0001100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001100001";
            uut_rst <= '0';
          WHEN "0001100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001100010";
            uut_rst <= '0';
          WHEN "0001100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001100011";
            uut_rst <= '0';
          WHEN "0001100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001100100";
            uut_rst <= '0';
          WHEN "0001100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001100101";
            uut_rst <= '0';
          WHEN "0001100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001100110";
            uut_rst <= '0';
          WHEN "0001100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001100111";
            uut_rst <= '0';
          WHEN "0001100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001101000";
            uut_rst <= '0';
          WHEN "0001101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001101001";
            uut_rst <= '0';
          WHEN "0001101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001101010";
            uut_rst <= '0';
          WHEN "0001101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001101011";
            uut_rst <= '0';
          WHEN "0001101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001101100";
            uut_rst <= '0';
          WHEN "0001101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001101101";
            uut_rst <= '0';
          WHEN "0001101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001101110";
            uut_rst <= '0';
          WHEN "0001101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001101111";
            uut_rst <= '0';
          WHEN "0001101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001110000";
            uut_rst <= '0';
          WHEN "0001110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001110001";
            uut_rst <= '0';
          WHEN "0001110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001110010";
            uut_rst <= '0';
          WHEN "0001110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001110011";
            uut_rst <= '0';
          WHEN "0001110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001110100";
            uut_rst <= '0';
          WHEN "0001110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001110101";
            uut_rst <= '0';
          WHEN "0001110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001110110";
            uut_rst <= '0';
          WHEN "0001110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001110111";
            uut_rst <= '0';
          WHEN "0001110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001111000";
            uut_rst <= '0';
          WHEN "0001111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001111001";
            uut_rst <= '0';
          WHEN "0001111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001111010";
            uut_rst <= '0';
          WHEN "0001111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001111011";
            uut_rst <= '0';
          WHEN "0001111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001111100";
            uut_rst <= '0';
          WHEN "0001111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001111101";
            uut_rst <= '0';
          WHEN "0001111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001111110";
            uut_rst <= '0';
          WHEN "0001111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0001111111";
            uut_rst <= '0';
          WHEN "0001111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010000000";
            uut_rst <= '0';
          WHEN "0010000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010000001";
            uut_rst <= '0';
          WHEN "0010000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010000010";
            uut_rst <= '0';
          WHEN "0010000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010000011";
            uut_rst <= '0';
          WHEN "0010000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010000100";
            uut_rst <= '0';
          WHEN "0010000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010000101";
            uut_rst <= '0';
          WHEN "0010000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010000110";
            uut_rst <= '0';
          WHEN "0010000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010000111";
            uut_rst <= '0';
          WHEN "0010000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010001000";
            uut_rst <= '0';
          WHEN "0010001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010001001";
            uut_rst <= '0';
          WHEN "0010001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010001010";
            uut_rst <= '0';
          WHEN "0010001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010001011";
            uut_rst <= '0';
          WHEN "0010001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010001100";
            uut_rst <= '0';
          WHEN "0010001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010001101";
            uut_rst <= '0';
          WHEN "0010001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010001110";
            uut_rst <= '0';
          WHEN "0010001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010001111";
            uut_rst <= '0';
          WHEN "0010001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010010000";
            uut_rst <= '0';
          WHEN "0010010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010010001";
            uut_rst <= '0';
          WHEN "0010010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010010010";
            uut_rst <= '0';
          WHEN "0010010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010010011";
            uut_rst <= '0';
          WHEN "0010010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010010100";
            uut_rst <= '0';
          WHEN "0010010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010010101";
            uut_rst <= '0';
          WHEN "0010010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010010110";
            uut_rst <= '0';
          WHEN "0010010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010010111";
            uut_rst <= '0';
          WHEN "0010010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010011000";
            uut_rst <= '0';
          WHEN "0010011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010011001";
            uut_rst <= '0';
          WHEN "0010011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010011010";
            uut_rst <= '0';
          WHEN "0010011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010011011";
            uut_rst <= '0';
          WHEN "0010011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010011100";
            uut_rst <= '0';
          WHEN "0010011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010011101";
            uut_rst <= '0';
          WHEN "0010011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010011110";
            uut_rst <= '0';
          WHEN "0010011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010011111";
            uut_rst <= '0';
          WHEN "0010011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010100000";
            uut_rst <= '0';
          WHEN "0010100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010100001";
            uut_rst <= '0';
          WHEN "0010100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010100010";
            uut_rst <= '0';
          WHEN "0010100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010100011";
            uut_rst <= '0';
          WHEN "0010100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010100100";
            uut_rst <= '0';
          WHEN "0010100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010100101";
            uut_rst <= '0';
          WHEN "0010100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010100110";
            uut_rst <= '0';
          WHEN "0010100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010100111";
            uut_rst <= '0';
          WHEN "0010100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010101000";
            uut_rst <= '0';
          WHEN "0010101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010101001";
            uut_rst <= '0';
          WHEN "0010101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010101010";
            uut_rst <= '0';
          WHEN "0010101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010101011";
            uut_rst <= '0';
          WHEN "0010101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010101100";
            uut_rst <= '0';
          WHEN "0010101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010101101";
            uut_rst <= '0';
          WHEN "0010101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010101110";
            uut_rst <= '0';
          WHEN "0010101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010101111";
            uut_rst <= '0';
          WHEN "0010101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010110000";
            uut_rst <= '0';
          WHEN "0010110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010110001";
            uut_rst <= '0';
          WHEN "0010110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010110010";
            uut_rst <= '0';
          WHEN "0010110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010110011";
            uut_rst <= '0';
          WHEN "0010110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010110100";
            uut_rst <= '0';
          WHEN "0010110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010110101";
            uut_rst <= '0';
          WHEN "0010110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010110110";
            uut_rst <= '0';
          WHEN "0010110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010110111";
            uut_rst <= '0';
          WHEN "0010110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010111000";
            uut_rst <= '0';
          WHEN "0010111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010111001";
            uut_rst <= '0';
          WHEN "0010111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010111010";
            uut_rst <= '0';
          WHEN "0010111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010111011";
            uut_rst <= '0';
          WHEN "0010111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010111100";
            uut_rst <= '0';
          WHEN "0010111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010111101";
            uut_rst <= '0';
          WHEN "0010111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010111110";
            uut_rst <= '0';
          WHEN "0010111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0010111111";
            uut_rst <= '0';
          WHEN "0010111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011000000";
            uut_rst <= '0';
          WHEN "0011000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011000001";
            uut_rst <= '0';
          WHEN "0011000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011000010";
            uut_rst <= '0';
          WHEN "0011000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011000011";
            uut_rst <= '0';
          WHEN "0011000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011000100";
            uut_rst <= '0';
          WHEN "0011000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011000101";
            uut_rst <= '0';
          WHEN "0011000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011000110";
            uut_rst <= '0';
          WHEN "0011000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011000111";
            uut_rst <= '0';
          WHEN "0011000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011001000";
            uut_rst <= '0';
          WHEN "0011001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011001001";
            uut_rst <= '0';
          WHEN "0011001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011001010";
            uut_rst <= '0';
          WHEN "0011001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011001011";
            uut_rst <= '0';
          WHEN "0011001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011001100";
            uut_rst <= '0';
          WHEN "0011001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011001101";
            uut_rst <= '0';
          WHEN "0011001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011001110";
            uut_rst <= '0';
          WHEN "0011001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011001111";
            uut_rst <= '0';
          WHEN "0011001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011010000";
            uut_rst <= '0';
          WHEN "0011010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011010001";
            uut_rst <= '0';
          WHEN "0011010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011010010";
            uut_rst <= '0';
          WHEN "0011010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011010011";
            uut_rst <= '0';
          WHEN "0011010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011010100";
            uut_rst <= '0';
          WHEN "0011010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011010101";
            uut_rst <= '0';
          WHEN "0011010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011010110";
            uut_rst <= '0';
          WHEN "0011010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011010111";
            uut_rst <= '0';
          WHEN "0011010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011011000";
            uut_rst <= '0';
          WHEN "0011011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011011001";
            uut_rst <= '0';
          WHEN "0011011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011011010";
            uut_rst <= '0';
          WHEN "0011011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011011011";
            uut_rst <= '0';
          WHEN "0011011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011011100";
            uut_rst <= '0';
          WHEN "0011011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011011101";
            uut_rst <= '0';
          WHEN "0011011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011011110";
            uut_rst <= '0';
          WHEN "0011011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011011111";
            uut_rst <= '0';
          WHEN "0011011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011100000";
            uut_rst <= '0';
          WHEN "0011100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011100001";
            uut_rst <= '0';
          WHEN "0011100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011100010";
            uut_rst <= '0';
          WHEN "0011100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011100011";
            uut_rst <= '0';
          WHEN "0011100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011100100";
            uut_rst <= '0';
          WHEN "0011100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011100101";
            uut_rst <= '0';
          WHEN "0011100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011100110";
            uut_rst <= '0';
          WHEN "0011100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011100111";
            uut_rst <= '0';
          WHEN "0011100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011101000";
            uut_rst <= '0';
          WHEN "0011101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011101001";
            uut_rst <= '0';
          WHEN "0011101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011101010";
            uut_rst <= '0';
          WHEN "0011101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011101011";
            uut_rst <= '0';
          WHEN "0011101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011101100";
            uut_rst <= '0';
          WHEN "0011101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011101101";
            uut_rst <= '0';
          WHEN "0011101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011101110";
            uut_rst <= '0';
          WHEN "0011101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011101111";
            uut_rst <= '0';
          WHEN "0011101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011110000";
            uut_rst <= '0';
          WHEN "0011110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011110001";
            uut_rst <= '0';
          WHEN "0011110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011110010";
            uut_rst <= '0';
          WHEN "0011110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011110011";
            uut_rst <= '0';
          WHEN "0011110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011110100";
            uut_rst <= '0';
          WHEN "0011110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011110101";
            uut_rst <= '0';
          WHEN "0011110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011110110";
            uut_rst <= '0';
          WHEN "0011110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011110111";
            uut_rst <= '0';
          WHEN "0011110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011111000";
            uut_rst <= '0';
          WHEN "0011111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011111001";
            uut_rst <= '0';
          WHEN "0011111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011111010";
            uut_rst <= '0';
          WHEN "0011111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011111011";
            uut_rst <= '0';
          WHEN "0011111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011111100";
            uut_rst <= '0';
          WHEN "0011111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011111101";
            uut_rst <= '0';
          WHEN "0011111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011111110";
            uut_rst <= '0';
          WHEN "0011111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0011111111";
            uut_rst <= '0';
          WHEN "0011111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100000000";
            uut_rst <= '0';
          WHEN "0100000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100000001";
            uut_rst <= '0';
          WHEN "0100000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100000010";
            uut_rst <= '0';
          WHEN "0100000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100000011";
            uut_rst <= '0';
          WHEN "0100000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100000100";
            uut_rst <= '0';
          WHEN "0100000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100000101";
            uut_rst <= '0';
          WHEN "0100000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100000110";
            uut_rst <= '0';
          WHEN "0100000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100000111";
            uut_rst <= '0';
          WHEN "0100000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100001000";
            uut_rst <= '0';
          WHEN "0100001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100001001";
            uut_rst <= '0';
          WHEN "0100001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100001010";
            uut_rst <= '0';
          WHEN "0100001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100001011";
            uut_rst <= '0';
          WHEN "0100001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100001100";
            uut_rst <= '0';
          WHEN "0100001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100001101";
            uut_rst <= '0';
          WHEN "0100001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100001110";
            uut_rst <= '0';
          WHEN "0100001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100001111";
            uut_rst <= '0';
          WHEN "0100001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100010000";
            uut_rst <= '0';
          WHEN "0100010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100010001";
            uut_rst <= '0';
          WHEN "0100010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100010010";
            uut_rst <= '0';
          WHEN "0100010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100010011";
            uut_rst <= '0';
          WHEN "0100010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100010100";
            uut_rst <= '0';
          WHEN "0100010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100010101";
            uut_rst <= '0';
          WHEN "0100010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100010110";
            uut_rst <= '0';
          WHEN "0100010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100010111";
            uut_rst <= '0';
          WHEN "0100010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100011000";
            uut_rst <= '0';
          WHEN "0100011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100011001";
            uut_rst <= '0';
          WHEN "0100011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100011010";
            uut_rst <= '0';
          WHEN "0100011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100011011";
            uut_rst <= '0';
          WHEN "0100011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100011100";
            uut_rst <= '0';
          WHEN "0100011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100011101";
            uut_rst <= '0';
          WHEN "0100011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100011110";
            uut_rst <= '0';
          WHEN "0100011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100011111";
            uut_rst <= '0';
          WHEN "0100011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100100000";
            uut_rst <= '0';
          WHEN "0100100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100100001";
            uut_rst <= '0';
          WHEN "0100100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100100010";
            uut_rst <= '0';
          WHEN "0100100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100100011";
            uut_rst <= '0';
          WHEN "0100100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100100100";
            uut_rst <= '0';
          WHEN "0100100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100100101";
            uut_rst <= '0';
          WHEN "0100100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100100110";
            uut_rst <= '0';
          WHEN "0100100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100100111";
            uut_rst <= '0';
          WHEN "0100100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100101000";
            uut_rst <= '0';
          WHEN "0100101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100101001";
            uut_rst <= '0';
          WHEN "0100101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100101010";
            uut_rst <= '0';
          WHEN "0100101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100101011";
            uut_rst <= '0';
          WHEN "0100101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100101100";
            uut_rst <= '0';
          WHEN "0100101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100101101";
            uut_rst <= '0';
          WHEN "0100101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100101110";
            uut_rst <= '0';
          WHEN "0100101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100101111";
            uut_rst <= '0';
          WHEN "0100101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100110000";
            uut_rst <= '0';
          WHEN "0100110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100110001";
            uut_rst <= '0';
          WHEN "0100110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100110010";
            uut_rst <= '0';
          WHEN "0100110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100110011";
            uut_rst <= '0';
          WHEN "0100110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100110100";
            uut_rst <= '0';
          WHEN "0100110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100110101";
            uut_rst <= '0';
          WHEN "0100110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100110110";
            uut_rst <= '0';
          WHEN "0100110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100110111";
            uut_rst <= '0';
          WHEN "0100110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100111000";
            uut_rst <= '0';
          WHEN "0100111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100111001";
            uut_rst <= '0';
          WHEN "0100111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100111010";
            uut_rst <= '0';
          WHEN "0100111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100111011";
            uut_rst <= '0';
          WHEN "0100111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100111100";
            uut_rst <= '0';
          WHEN "0100111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100111101";
            uut_rst <= '0';
          WHEN "0100111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100111110";
            uut_rst <= '0';
          WHEN "0100111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0100111111";
            uut_rst <= '0';
          WHEN "0100111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101000000";
            uut_rst <= '0';
          WHEN "0101000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101000001";
            uut_rst <= '0';
          WHEN "0101000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101000010";
            uut_rst <= '0';
          WHEN "0101000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101000011";
            uut_rst <= '0';
          WHEN "0101000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101000100";
            uut_rst <= '0';
          WHEN "0101000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101000101";
            uut_rst <= '0';
          WHEN "0101000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101000110";
            uut_rst <= '0';
          WHEN "0101000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101000111";
            uut_rst <= '0';
          WHEN "0101000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101001000";
            uut_rst <= '0';
          WHEN "0101001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101001001";
            uut_rst <= '0';
          WHEN "0101001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101001010";
            uut_rst <= '0';
          WHEN "0101001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101001011";
            uut_rst <= '0';
          WHEN "0101001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101001100";
            uut_rst <= '0';
          WHEN "0101001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101001101";
            uut_rst <= '0';
          WHEN "0101001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101001110";
            uut_rst <= '0';
          WHEN "0101001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101001111";
            uut_rst <= '0';
          WHEN "0101001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101010000";
            uut_rst <= '0';
          WHEN "0101010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101010001";
            uut_rst <= '0';
          WHEN "0101010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101010010";
            uut_rst <= '0';
          WHEN "0101010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101010011";
            uut_rst <= '0';
          WHEN "0101010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101010100";
            uut_rst <= '0';
          WHEN "0101010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101010101";
            uut_rst <= '0';
          WHEN "0101010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101010110";
            uut_rst <= '0';
          WHEN "0101010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101010111";
            uut_rst <= '0';
          WHEN "0101010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101011000";
            uut_rst <= '0';
          WHEN "0101011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101011001";
            uut_rst <= '0';
          WHEN "0101011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101011010";
            uut_rst <= '0';
          WHEN "0101011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101011011";
            uut_rst <= '0';
          WHEN "0101011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101011100";
            uut_rst <= '0';
          WHEN "0101011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101011101";
            uut_rst <= '0';
          WHEN "0101011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101011110";
            uut_rst <= '0';
          WHEN "0101011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101011111";
            uut_rst <= '0';
          WHEN "0101011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101100000";
            uut_rst <= '0';
          WHEN "0101100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101100001";
            uut_rst <= '0';
          WHEN "0101100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101100010";
            uut_rst <= '0';
          WHEN "0101100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101100011";
            uut_rst <= '0';
          WHEN "0101100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101100100";
            uut_rst <= '0';
          WHEN "0101100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101100101";
            uut_rst <= '0';
          WHEN "0101100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101100110";
            uut_rst <= '0';
          WHEN "0101100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101100111";
            uut_rst <= '0';
          WHEN "0101100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101101000";
            uut_rst <= '0';
          WHEN "0101101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101101001";
            uut_rst <= '0';
          WHEN "0101101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101101010";
            uut_rst <= '0';
          WHEN "0101101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101101011";
            uut_rst <= '0';
          WHEN "0101101011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101101100";
            uut_rst <= '0';
          WHEN "0101101100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101101101";
            uut_rst <= '0';
          WHEN "0101101101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101101110";
            uut_rst <= '0';
          WHEN "0101101110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101101111";
            uut_rst <= '0';
          WHEN "0101101111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101110000";
            uut_rst <= '0';
          WHEN "0101110000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101110001";
            uut_rst <= '0';
          WHEN "0101110001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101110010";
            uut_rst <= '0';
          WHEN "0101110010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101110011";
            uut_rst <= '0';
          WHEN "0101110011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101110100";
            uut_rst <= '0';
          WHEN "0101110100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101110101";
            uut_rst <= '0';
          WHEN "0101110101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101110110";
            uut_rst <= '0';
          WHEN "0101110110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101110111";
            uut_rst <= '0';
          WHEN "0101110111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101111000";
            uut_rst <= '0';
          WHEN "0101111000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101111001";
            uut_rst <= '0';
          WHEN "0101111001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101111010";
            uut_rst <= '0';
          WHEN "0101111010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101111011";
            uut_rst <= '0';
          WHEN "0101111011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101111100";
            uut_rst <= '0';
          WHEN "0101111100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101111101";
            uut_rst <= '0';
          WHEN "0101111101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101111110";
            uut_rst <= '0';
          WHEN "0101111110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0101111111";
            uut_rst <= '0';
          WHEN "0101111111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110000000";
            uut_rst <= '0';
          WHEN "0110000000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110000001";
            uut_rst <= '0';
          WHEN "0110000001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110000010";
            uut_rst <= '0';
          WHEN "0110000010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110000011";
            uut_rst <= '0';
          WHEN "0110000011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110000100";
            uut_rst <= '0';
          WHEN "0110000100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110000101";
            uut_rst <= '0';
          WHEN "0110000101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110000110";
            uut_rst <= '0';
          WHEN "0110000110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110000111";
            uut_rst <= '0';
          WHEN "0110000111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110001000";
            uut_rst <= '0';
          WHEN "0110001000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110001001";
            uut_rst <= '0';
          WHEN "0110001001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110001010";
            uut_rst <= '0';
          WHEN "0110001010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110001011";
            uut_rst <= '0';
          WHEN "0110001011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110001100";
            uut_rst <= '0';
          WHEN "0110001100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110001101";
            uut_rst <= '0';
          WHEN "0110001101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110001110";
            uut_rst <= '0';
          WHEN "0110001110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110001111";
            uut_rst <= '0';
          WHEN "0110001111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110010000";
            uut_rst <= '0';
          WHEN "0110010000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110010001";
            uut_rst <= '0';
          WHEN "0110010001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110010010";
            uut_rst <= '0';
          WHEN "0110010010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110010011";
            uut_rst <= '0';
          WHEN "0110010011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110010100";
            uut_rst <= '0';
          WHEN "0110010100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110010101";
            uut_rst <= '0';
          WHEN "0110010101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110010110";
            uut_rst <= '0';
          WHEN "0110010110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110010111";
            uut_rst <= '0';
          WHEN "0110010111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110011000";
            uut_rst <= '0';
          WHEN "0110011000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110011001";
            uut_rst <= '0';
          WHEN "0110011001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110011010";
            uut_rst <= '0';
          WHEN "0110011010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110011011";
            uut_rst <= '0';
          WHEN "0110011011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110011100";
            uut_rst <= '0';
          WHEN "0110011100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110011101";
            uut_rst <= '0';
          WHEN "0110011101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110011110";
            uut_rst <= '0';
          WHEN "0110011110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110011111";
            uut_rst <= '0';
          WHEN "0110011111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110100000";
            uut_rst <= '0';
          WHEN "0110100000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110100001";
            uut_rst <= '0';
          WHEN "0110100001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110100010";
            uut_rst <= '0';
          WHEN "0110100010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110100011";
            uut_rst <= '0';
          WHEN "0110100011" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110100100";
            uut_rst <= '0';
          WHEN "0110100100" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110100101";
            uut_rst <= '0';
          WHEN "0110100101" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110100110";
            uut_rst <= '0';
          WHEN "0110100110" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110100111";
            uut_rst <= '0';
          WHEN "0110100111" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110101000";
            uut_rst <= '0';
          WHEN "0110101000" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110101001";
            uut_rst <= '0';
          WHEN "0110101001" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110101010";
            uut_rst <= '0';
          WHEN "0110101010" =>
            uut_input_load <= '0';
            uut_a_0_0 <= "000000000000000000000000000";
            uut_a_0_1 <= "000000000000000000000000000";
            uut_a_0_2 <= "000000000000000000000000000";
            uut_a_0_3 <= "000000000000000000000000000";
            uut_a_0_4 <= "000000000000000000000000000";
            uut_a_0_5 <= "000000000000000000000000000";
            uut_a_1_0 <= "000000000000000000000000000";
            uut_a_1_1 <= "000000000000000000000000000";
            uut_a_1_2 <= "000000000000000000000000000";
            uut_a_1_3 <= "000000000000000000000000000";
            uut_a_1_4 <= "000000000000000000000000000";
            uut_a_1_5 <= "000000000000000000000000000";
            uut_a_2_0 <= "000000000000000000000000000";
            uut_a_2_1 <= "000000000000000000000000000";
            uut_a_2_2 <= "000000000000000000000000000";
            uut_a_2_3 <= "000000000000000000000000000";
            uut_a_2_4 <= "000000000000000000000000000";
            uut_a_2_5 <= "000000000000000000000000000";
            uut_a_3_0 <= "000000000000000000000000000";
            uut_a_3_1 <= "000000000000000000000000000";
            uut_a_3_2 <= "000000000000000000000000000";
            uut_a_3_3 <= "000000000000000000000000000";
            uut_a_3_4 <= "000000000000000000000000000";
            uut_a_3_5 <= "000000000000000000000000000";
            uut_a_4_0 <= "000000000000000000000000000";
            uut_a_4_1 <= "000000000000000000000000000";
            uut_a_4_2 <= "000000000000000000000000000";
            uut_a_4_3 <= "000000000000000000000000000";
            uut_a_4_4 <= "000000000000000000000000000";
            uut_a_4_5 <= "000000000000000000000000000";
            uut_a_5_0 <= "000000000000000000000000000";
            uut_a_5_1 <= "000000000000000000000000000";
            uut_a_5_2 <= "000000000000000000000000000";
            uut_a_5_3 <= "000000000000000000000000000";
            uut_a_5_4 <= "000000000000000000000000000";
            uut_a_5_5 <= "000000000000000000000000000";
            uut_b_0 <= "000000000000000000000000000";
            uut_b_1 <= "000000000000000000000000000";
            uut_b_2 <= "000000000000000000000000000";
            uut_b_3 <= "000000000000000000000000000";
            uut_b_4 <= "000000000000000000000000000";
            uut_b_5 <= "000000000000000000000000000";
            state <= "0110101011";
            uut_rst <= '0';
          WHEN "0110101011" =>
            state <= "0110101100";
            uut_rst <= '0';
          WHEN "0110101100" =>
            state <= "0110101101";
            uut_rst <= '0';
          WHEN "0110101101" =>
            state <= "0110101110";
            uut_rst <= '0';
          WHEN "0110101110" =>
            state <= "0110101111";
            uut_rst <= '0';
          WHEN "0110101111" =>
            state <= "0110110000";
            uut_rst <= '0';
          WHEN "0110110000" =>
            state <= "0110110001";
            uut_rst <= '0';
          WHEN "0110110001" =>
            state <= "0110110010";
            uut_rst <= '0';
          WHEN "0110110010" =>
            state <= "0110110011";
            uut_rst <= '0';
          WHEN "0110110011" =>
            state <= "0110110100";
            uut_rst <= '0';
          WHEN "0110110100" =>
            state <= "0110110101";
            uut_rst <= '0';
          WHEN "0110110101" =>
            state <= "0110110110";
            uut_rst <= '0';
          WHEN "0110110110" =>
            state <= "0110110111";
            uut_rst <= '0';
          WHEN "0110110111" =>
            state <= "0110111000";
            uut_rst <= '0';
          WHEN "0110111000" =>
            state <= "0110111001";
            uut_rst <= '0';
          WHEN "0110111001" =>
            state <= "0110111010";
            uut_rst <= '0';
          WHEN "0110111010" =>
            state <= "0110111011";
            uut_rst <= '0';
          WHEN "0110111011" =>
            state <= "0110111100";
            uut_rst <= '0';
          WHEN "0110111100" =>
            state <= "0110111101";
            uut_rst <= '0';
          WHEN "0110111101" =>
            state <= "0110111110";
            uut_rst <= '0';
          WHEN "0110111110" =>
            state <= "0110111111";
            uut_rst <= '0';
          WHEN "0110111111" =>
            state <= "0111000000";
            uut_rst <= '0';
          WHEN "0111000000" =>
            state <= "0111000001";
            uut_rst <= '0';
          WHEN "0111000001" =>
            state <= "0111000010";
            uut_rst <= '0';
          WHEN "0111000010" =>
            state <= "0111000011";
            uut_rst <= '0';
          WHEN "0111000011" =>
            state <= "0111000100";
            uut_rst <= '0';
          WHEN "0111000100" =>
            state <= "0111000101";
            uut_rst <= '0';
          WHEN "0111000101" =>
            state <= "0111000110";
            uut_rst <= '0';
          WHEN "0111000110" =>
            state <= "0111000111";
            uut_rst <= '0';
          WHEN "0111000111" =>
            state <= "0111001000";
            uut_rst <= '0';
          WHEN "0111001000" =>
            state <= "0111001001";
            uut_rst <= '0';
          WHEN "0111001001" =>
            state <= "0111001010";
            uut_rst <= '0';
          WHEN "0111001010" =>
            state <= "0111001011";
            uut_rst <= '0';
          WHEN "0111001011" =>
            state <= "0111001100";
            uut_rst <= '0';
          WHEN "0111001100" =>
            state <= "0111001101";
            uut_rst <= '0';
          WHEN "0111001101" =>
            state <= "0111001110";
            uut_rst <= '0';
          WHEN "0111001110" =>
            state <= "0111001111";
            uut_rst <= '0';
          WHEN "0111001111" =>
            state <= "0111010000";
            uut_rst <= '0';
          WHEN "0111010000" =>
            state <= "0111010001";
            uut_rst <= '0';
          WHEN "0111010001" =>
            state <= "0111010010";
            uut_rst <= '0';
          WHEN "0111010010" =>
            state <= "0111010011";
            uut_rst <= '0';
          WHEN "0111010011" =>
            state <= "0111010100";
            uut_rst <= '0';
          WHEN "0111010100" =>
            state <= "0111010101";
            uut_rst <= '0';
          WHEN "0111010101" =>
            state <= "0111010110";
            uut_rst <= '0';
          WHEN "0111010110" =>
            state <= "0111010111";
            uut_rst <= '0';
          WHEN "0111010111" =>
            state <= "0111011000";
            uut_rst <= '0';
          WHEN "0111011000" =>
            state <= "0111011001";
            uut_rst <= '0';
          WHEN "0111011001" =>
            state <= "0111011010";
            uut_rst <= '0';
          WHEN "0111011010" =>
            state <= "0111011011";
            uut_rst <= '0';
          WHEN "0111011011" =>
            state <= "0111011100";
            uut_rst <= '0';
          WHEN "0111011100" =>
            state <= "0111011101";
            uut_rst <= '0';
          WHEN "0111011101" =>
            state <= "0111011110";
            uut_rst <= '0';
          WHEN "0111011110" =>
            state <= "0111011111";
            uut_rst <= '0';
          WHEN "0111011111" =>
            state <= "0111100000";
            uut_rst <= '0';
          WHEN "0111100000" =>
            state <= "0111100001";
            uut_rst <= '0';
          WHEN "0111100001" =>
            state <= "0111100010";
            uut_rst <= '0';
          WHEN "0111100010" =>
            state <= "0111100011";
            uut_rst <= '0';
          WHEN "0111100011" =>
            state <= "0111100100";
            uut_rst <= '0';
          WHEN "0111100100" =>
            state <= "0111100101";
            uut_rst <= '0';
          WHEN "0111100101" =>
            state <= "0111100110";
            uut_rst <= '0';
          WHEN "0111100110" =>
            state <= "0111100111";
            uut_rst <= '0';
          WHEN "0111100111" =>
            state <= "0111101000";
            uut_rst <= '0';
          WHEN "0111101000" =>
            state <= "0111101001";
            uut_rst <= '0';
          WHEN "0111101001" =>
            state <= "0111101010";
            uut_rst <= '0';
          WHEN "0111101010" =>
            state <= "0111101011";
            uut_rst <= '0';
          WHEN "0111101011" =>
            state <= "0111101100";
            uut_rst <= '0';
          WHEN "0111101100" =>
            state <= "0111101101";
            uut_rst <= '0';
          WHEN "0111101101" =>
            state <= "0111101110";
            uut_rst <= '0';
          WHEN "0111101110" =>
            state <= "0111101111";
            uut_rst <= '0';
          WHEN "0111101111" =>
            state <= "0111110000";
            uut_rst <= '0';
          WHEN "0111110000" =>
            state <= "0111110001";
            uut_rst <= '0';
          WHEN "0111110001" =>
            state <= "0111110010";
            uut_rst <= '0';
          WHEN "0111110010" =>
            state <= "0111110011";
            uut_rst <= '0';
          WHEN "0111110011" =>
            state <= "0111110100";
            uut_rst <= '0';
          WHEN "0111110100" =>
            state <= "0111110101";
            uut_rst <= '0';
          WHEN "0111110101" =>
            state <= "0111110110";
            uut_rst <= '0';
          WHEN "0111110110" =>
            state <= "0111110111";
            uut_rst <= '0';
          WHEN "0111110111" =>
            state <= "0111111000";
            uut_rst <= '0';
          WHEN "0111111000" =>
            state <= "0111111001";
            uut_rst <= '0';
          WHEN "0111111001" =>
            state <= "0111111010";
            uut_rst <= '0';
          WHEN "0111111010" =>
            state <= "0111111011";
            uut_rst <= '0';
          WHEN "0111111011" =>
            state <= "0111111100";
            uut_rst <= '0';
          WHEN "0111111100" =>
            state <= "0111111101";
            uut_rst <= '0';
          WHEN "0111111101" =>
            state <= "0111111110";
            uut_rst <= '0';
          WHEN "0111111110" =>
            state <= "0111111111";
            uut_rst <= '0';
          WHEN "0111111111" =>
            state <= "1000000000";
            uut_rst <= '0';
          WHEN "1000000000" =>
            state <= "1000000001";
            uut_rst <= '0';
          WHEN "1000000001" =>
            state <= "1000000010";
            uut_rst <= '0';
          WHEN "1000000010" =>
            state <= "1000000011";
            uut_rst <= '0';
          WHEN "1000000011" =>
            state <= "1000000100";
            uut_rst <= '0';
          WHEN "1000000100" =>
            state <= "1000000101";
            uut_rst <= '0';
          WHEN "1000000101" =>
            state <= "1000000110";
            uut_rst <= '0';
          WHEN "1000000110" =>
            state <= "1000000111";
            uut_rst <= '0';
          WHEN "1000000111" =>
            state <= "1000001000";
            uut_rst <= '0';
          WHEN "1000001000" =>
            state <= "1000001001";
            uut_rst <= '0';
          WHEN "1000001001" =>
            state <= "1000001010";
            uut_rst <= '0';
          WHEN "1000001010" =>
            state <= "1000001011";
            uut_rst <= '0';
          WHEN "1000001011" =>
            state <= "1000001100";
            uut_rst <= '0';
          WHEN "1000001100" =>
            state <= "1000001101";
            uut_rst <= '0';
          WHEN "1000001101" =>
            state <= "1000001110";
            uut_rst <= '0';
          WHEN "1000001110" =>
            state <= "1000001111";
            uut_rst <= '0';
          WHEN "1000001111" =>
            state <= "1000010000";
            uut_rst <= '0';
          WHEN "1000010000" =>
            state <= "1000010001";
            uut_rst <= '0';
          WHEN "1000010001" =>
            state <= "1000010010";
            uut_rst <= '0';
          WHEN "1000010010" =>
            state <= "1000010011";
            uut_rst <= '0';
          WHEN "1000010011" =>
            state <= "1000010100";
            uut_rst <= '0';
          WHEN "1000010100" =>
            state <= "1000010101";
            uut_rst <= '0';
          WHEN "1000010101" =>
            state <= "1000010110";
            uut_rst <= '0';
          WHEN "1000010110" =>
            state <= "1000010111";
            uut_rst <= '0';
          WHEN "1000010111" =>
            state <= "1000011000";
            uut_rst <= '0';
          WHEN "1000011000" =>
            state <= "1000011001";
            uut_rst <= '0';
          WHEN "1000011001" =>
            state <= "1000011010";
            uut_rst <= '0';
          WHEN "1000011010" =>
            state <= "1000011011";
            uut_rst <= '0';
          WHEN "1000011011" =>
            state <= "1000011100";
            uut_rst <= '0';
          WHEN "1000011100" =>
            state <= "1000011101";
            uut_rst <= '0';
          WHEN "1000011101" =>
            state <= "1000011110";
            uut_rst <= '0';
          WHEN "1000011110" =>
            state <= "1000011111";
            uut_rst <= '0';
          WHEN "1000011111" =>
            state <= "1000100000";
            uut_rst <= '0';
          WHEN "1000100000" =>
            state <= "1000100001";
            uut_rst <= '0';
          WHEN "1000100001" =>
            state <= "1000100010";
            uut_rst <= '0';
          WHEN "1000100010" =>
            state <= "1000100011";
            uut_rst <= '0';
          WHEN "1000100011" =>
            state <= "1000100100";
            uut_rst <= '0';
          WHEN "1000100100" =>
            state <= "1000100101";
            uut_rst <= '0';
          WHEN "1000100101" =>
            state <= "1000100110";
            uut_rst <= '0';
          WHEN "1000100110" =>
            state <= "1000100111";
            uut_rst <= '0';
          WHEN "1000100111" =>
            state <= "1000101000";
            uut_rst <= '0';
          WHEN "1000101000" =>
            state <= "1000101001";
            uut_rst <= '0';
          WHEN "1000101001" =>
            state <= "1000101010";
            uut_rst <= '0';
          WHEN "1000101010" =>
            state <= "1000101011";
            uut_rst <= '0';
          WHEN "1000101011" =>
            state <= "1000101100";
            uut_rst <= '0';
          WHEN "1000101100" =>
            state <= "1000101101";
            uut_rst <= '0';
          WHEN "1000101101" =>
            state <= "1000101110";
            uut_rst <= '0';
          WHEN "1000101110" =>
            state <= "1000101111";
            uut_rst <= '0';
          WHEN "1000101111" =>
            state <= "1000110000";
            uut_rst <= '0';
          WHEN "1000110000" =>
            state <= "1000110001";
            uut_rst <= '0';
          WHEN "1000110001" =>
            state <= "1000110010";
            uut_rst <= '0';
          WHEN "1000110010" =>
            state <= "1000110011";
            uut_rst <= '0';
          WHEN "1000110011" =>
            state <= "1000110100";
            uut_rst <= '0';
          WHEN "1000110100" =>
            state <= "1000110101";
            uut_rst <= '0';
          WHEN "1000110101" =>
            state <= "1000110110";
            uut_rst <= '0';
          WHEN "1000110110" =>
            state <= "1000110111";
            uut_rst <= '0';
          WHEN "1000110111" =>
            state <= "1000111000";
            uut_rst <= '0';
          WHEN "1000111000" =>
            state <= "1000111001";
            uut_rst <= '0';
          WHEN "1000111001" =>
            state <= "1000111010";
            uut_rst <= '0';
          WHEN "1000111010" =>
            state <= "1000111011";
            uut_rst <= '0';
          WHEN "1000111011" =>
            state <= "1000111100";
            uut_rst <= '0';
          WHEN "1000111100" =>
            state <= "1000111101";
            uut_rst <= '0';
          WHEN "1000111101" =>
            state <= "1000111110";
            uut_rst <= '0';
          WHEN "1000111110" =>
            state <= "1000111111";
            uut_rst <= '0';
          WHEN "1000111111" =>
            state <= "1001000000";
            uut_rst <= '0';
          WHEN "1001000000" =>
            state <= "1001000001";
            uut_rst <= '0';
          WHEN "1001000001" =>
            state <= "1001000010";
            uut_rst <= '0';
          WHEN "1001000010" =>
            state <= "1001000011";
            uut_rst <= '0';
          WHEN "1001000011" =>
            state <= "1001000100";
            uut_rst <= '0';
          WHEN "1001000100" =>
            state <= "1001000101";
            uut_rst <= '0';
          WHEN "1001000101" =>
            state <= "1001000110";
            uut_rst <= '0';
          WHEN "1001000110" =>
            state <= "1001000111";
            uut_rst <= '0';
          WHEN "1001000111" =>
            state <= "1001001000";
            uut_rst <= '0';
          WHEN "1001001000" =>
            state <= "1001001001";
            uut_rst <= '0';
          WHEN "1001001001" =>
            state <= "1001001010";
            uut_rst <= '0';
          WHEN "1001001010" =>
            state <= "1001001011";
            uut_rst <= '0';
          WHEN "1001001011" =>
            state <= "1001001100";
            uut_rst <= '0';
          WHEN "1001001100" =>
            state <= "1001001101";
            uut_rst <= '0';
          WHEN "1001001101" =>
            state <= "1001001110";
            uut_rst <= '0';
          WHEN "1001001110" =>
            state <= "1001001111";
            uut_rst <= '0';
          WHEN "1001001111" =>
            state <= "1001010000";
            uut_rst <= '0';
          WHEN "1001010000" =>
            state <= "1001010001";
            uut_rst <= '0';
          WHEN "1001010001" =>
            state <= "1001010010";
            uut_rst <= '0';
          WHEN "1001010010" =>
            state <= "1001010011";
            uut_rst <= '0';
          WHEN "1001010011" =>
            state <= "1001010100";
            uut_rst <= '0';
          WHEN "1001010100" =>
            state <= "1001010101";
            uut_rst <= '0';
          WHEN "1001010101" =>
            state <= "1001010110";
            uut_rst <= '0';
          WHEN "1001010110" =>
            state <= "1001010111";
            uut_rst <= '0';
          WHEN "1001010111" =>
            state <= "1001011000";
            uut_rst <= '0';
          WHEN "1001011000" =>
            state <= "1001011001";
            uut_rst <= '0';
          WHEN "1001011001" =>
            state <= "1001011010";
            uut_rst <= '0';
          WHEN "1001011010" =>
            state <= "1001011011";
            uut_rst <= '0';
          WHEN "1001011011" =>
            state <= "1001011100";
            uut_rst <= '0';
          WHEN "1001011100" =>
            state <= "1001011101";
            uut_rst <= '0';
          WHEN "1001011101" =>
            state <= "1001011110";
            uut_rst <= '0';
          WHEN "1001011110" =>
            state <= "1001011111";
            uut_rst <= '0';
          WHEN "1001011111" =>
            state <= "1001100000";
            uut_rst <= '0';
          WHEN "1001100000" =>
            state <= "1001100001";
            uut_rst <= '0';
          WHEN "1001100001" =>
            state <= "1001100010";
            uut_rst <= '0';
          WHEN "1001100010" =>
            state <= "1001100011";
            uut_rst <= '0';
          WHEN "1001100011" =>
            state <= "1001100100";
            uut_rst <= '0';
          WHEN "1001100100" =>
            state <= "1001100101";
            uut_rst <= '0';
          WHEN "1001100101" =>
            state <= "1001100110";
            uut_rst <= '0';
          WHEN "1001100110" =>
            state <= "1001100111";
            uut_rst <= '0';
          WHEN "1001100111" =>
            state <= "1001101000";
            uut_rst <= '0';
          WHEN "1001101000" =>
            state <= "1001101001";
            uut_rst <= '0';
          WHEN "1001101001" =>
            state <= "1001101010";
            uut_rst <= '0';
          WHEN "1001101010" =>
            state <= "1001101011";
            uut_rst <= '0';
          WHEN "1001101011" =>
            state <= "1001101100";
            uut_rst <= '0';
          WHEN "1001101100" =>
            state <= "1001101101";
            uut_rst <= '0';
          WHEN "1001101101" =>
            state <= "1001101110";
            uut_rst <= '0';
          WHEN "1001101110" =>
            state <= "1001101111";
            uut_rst <= '0';
          WHEN "1001101111" =>
            state <= "1001110000";
            uut_rst <= '0';
          WHEN "1001110000" =>
            state <= "1001110001";
            uut_rst <= '0';
          WHEN "1001110001" =>
            state <= "1001110010";
            uut_rst <= '0';
          WHEN "1001110010" =>
            state <= "1001110011";
            uut_rst <= '0';
          WHEN "1001110011" =>
            state <= "1001110100";
            uut_rst <= '0';
          WHEN "1001110100" =>
            state <= "1001110101";
            uut_rst <= '0';
          WHEN "1001110101" =>
            state <= "1001110110";
            uut_rst <= '0';
          WHEN "1001110110" =>
            state <= "1001110111";
            uut_rst <= '0';
          WHEN "1001110111" =>
            state <= "1001111000";
            uut_rst <= '0';
          WHEN "1001111000" =>
            state <= "1001111001";
            uut_rst <= '0';
          WHEN "1001111001" =>
            state <= "1001111010";
            uut_rst <= '0';
          WHEN "1001111010" =>
            state <= "1001111011";
            uut_rst <= '0';
          WHEN "1001111011" =>
            state <= "1001111100";
            uut_rst <= '0';
          WHEN "1001111100" =>
            state <= "1001111101";
            uut_rst <= '0';
          WHEN "1001111101" =>
            state <= "1001111110";
            uut_rst <= '0';
          WHEN "1001111110" =>
            state <= "1001111111";
            uut_rst <= '0';
          WHEN "1001111111" =>
            state <= "1010000000";
            uut_rst <= '0';
          WHEN "1010000000" =>
            state <= "1010000001";
            uut_rst <= '0';
          WHEN "1010000001" =>
            state <= "1010000010";
            uut_rst <= '0';
          WHEN "1010000010" =>
            state <= "1010000011";
            uut_rst <= '0';
          WHEN "1010000011" =>
            state <= "1010000100";
            uut_rst <= '0';
          WHEN "1010000100" =>
            state <= "1010000101";
            uut_rst <= '0';
          WHEN "1010000101" =>
            state <= "1010000110";
            uut_rst <= '0';
          WHEN "1010000110" =>
            state <= "1010000111";
            uut_rst <= '0';
          WHEN "1010000111" =>
            state <= "1010001000";
            uut_rst <= '0';
          WHEN "1010001000" =>
            state <= "1010001001";
            uut_rst <= '0';
          WHEN "1010001001" =>
            state <= "1010001010";
            uut_rst <= '0';
          WHEN "1010001010" =>
            state <= "1010001011";
            uut_rst <= '0';
          WHEN "1010001011" =>
            state <= "1010001100";
            uut_rst <= '0';
          WHEN "1010001100" =>
            state <= "1010001101";
            uut_rst <= '0';
          WHEN "1010001101" =>
            state <= "1010001110";
            uut_rst <= '0';
          WHEN "1010001110" =>
            state <= "1010001111";
            uut_rst <= '0';
          WHEN "1010001111" =>
            state <= "1010010000";
            uut_rst <= '0';
          WHEN "1010010000" =>
            state <= "1010010001";
            uut_rst <= '0';
          WHEN "1010010001" =>
            state <= "1010010010";
            uut_rst <= '0';
          WHEN "1010010010" =>
            state <= "1010010011";
            uut_rst <= '0';
          WHEN "1010010011" =>
            state <= "1010010100";
            uut_rst <= '0';
          WHEN "1010010100" =>
            state <= "1010010101";
            uut_rst <= '0';
          WHEN "1010010101" =>
            state <= "1010010110";
            uut_rst <= '0';
          WHEN "1010010110" =>
            state <= "1010010111";
            uut_rst <= '0';
          WHEN "1010010111" =>
            state <= "1010011000";
            uut_rst <= '0';
          WHEN "1010011000" =>
            state <= "1010011001";
            uut_rst <= '0';
          WHEN "1010011001" =>
            state <= "1010011010";
            uut_rst <= '0';
          WHEN "1010011010" =>
            state <= "1010011011";
            uut_rst <= '0';
          WHEN "1010011011" =>
            state <= "1010011100";
            uut_rst <= '0';
          WHEN "1010011100" =>
            state <= "1010011101";
            uut_rst <= '0';
          WHEN "1010011101" =>
            state <= "1010011110";
            uut_rst <= '0';
          WHEN "1010011110" =>
            state <= "1010011111";
            uut_rst <= '0';
          WHEN "1010011111" =>
            state <= "1010100000";
            uut_rst <= '0';
          WHEN "1010100000" =>
            state <= "1010100001";
            uut_rst <= '0';
          WHEN "1010100001" =>
            state <= "1010100010";
            uut_rst <= '0';
          WHEN "1010100010" =>
            state <= "1010100011";
            uut_rst <= '0';
          WHEN "1010100011" =>
            state <= "1010100100";
            uut_rst <= '0';
          WHEN "1010100100" =>
            state <= "1010100101";
            uut_rst <= '0';
          WHEN "1010100101" =>
            state <= "1010100110";
            uut_rst <= '0';
          WHEN "1010100110" =>
            state <= "1010100111";
            uut_rst <= '0';
          WHEN "1010100111" =>
            state <= "1010101000";
            uut_rst <= '0';
          WHEN "1010101000" =>
            state <= "1010101001";
            uut_rst <= '0';
          WHEN "1010101001" =>
            state <= "1010101010";
            uut_rst <= '0';
          WHEN "1010101010" =>
            state <= "1010101011";
            uut_rst <= '0';
          WHEN "1010101011" =>
            state <= "1010101100";
            uut_rst <= '0';
          WHEN "1010101100" =>
            state <= "1010101101";
            uut_rst <= '0';
          WHEN "1010101101" =>
            state <= "1010101110";
            uut_rst <= '0';
          WHEN "1010101110" =>
            state <= "1010101111";
            uut_rst <= '0';
          WHEN "1010101111" =>
            state <= "1010110000";
            uut_rst <= '0';
          WHEN "1010110000" =>
            state <= "1010110001";
            uut_rst <= '0';
          WHEN "1010110001" =>
            state <= "1010110010";
            uut_rst <= '0';
          WHEN "1010110010" =>
            state <= "1010110011";
            uut_rst <= '0';
          WHEN "1010110011" =>
            state <= "1010110100";
            uut_rst <= '0';
          WHEN "1010110100" =>
            state <= "1010110101";
            uut_rst <= '0';
          WHEN "1010110101" =>
            state <= "1010110110";
            uut_rst <= '0';
          WHEN "1010110110" =>
            state <= "1010110111";
            uut_rst <= '0';
          WHEN "1010110111" =>
            state <= "1010111000";
            uut_rst <= '0';
          WHEN "1010111000" =>
            state <= "1010111001";
            uut_rst <= '0';
          WHEN "1010111001" =>
            state <= "1010111010";
            uut_rst <= '0';
          WHEN "1010111010" =>
            state <= "1010111011";
            uut_rst <= '0';
          WHEN "1010111011" =>
            state <= "1010111100";
            uut_rst <= '0';
          WHEN "1010111100" =>
            state <= "1010111101";
            uut_rst <= '0';
          WHEN "1010111101" =>
            state <= "1010111110";
            uut_rst <= '0';
          WHEN "1010111110" =>
            state <= "1010111111";
            uut_rst <= '0';
          WHEN "1010111111" =>
            state <= "1011000000";
            uut_rst <= '0';
          WHEN "1011000000" =>
            state <= "1011000001";
            uut_rst <= '0';
          WHEN "1011000001" =>
            state <= "1011000010";
            uut_rst <= '0';
          WHEN "1011000010" =>
            state <= "1011000011";
            uut_rst <= '0';
          WHEN "1011000011" =>
            state <= "1011000100";
            uut_rst <= '0';
          WHEN "1011000100" =>
            state <= "1011000101";
            uut_rst <= '0';
          WHEN "1011000101" =>
            state <= "1011000110";
            uut_rst <= '0';
          WHEN "1011000110" =>
            state <= "1011000111";
            uut_rst <= '0';
          WHEN "1011000111" =>
            state <= "1011001000";
            uut_rst <= '0';
          WHEN "1011001000" =>
            state <= "1011001001";
            uut_rst <= '0';
          WHEN "1011001001" =>
            state <= "1011001010";
            uut_rst <= '0';
          WHEN "1011001010" =>
            state <= "1011001011";
            uut_rst <= '0';
          WHEN "1011001011" =>
            state <= "1011001100";
            uut_rst <= '0';
          WHEN "1011001100" =>
            state <= "1011001101";
            uut_rst <= '0';
          WHEN "1011001101" =>
            state <= "1011001110";
            uut_rst <= '0';
          WHEN "1011001110" =>
            state <= "1011001111";
            uut_rst <= '0';
          WHEN "1011001111" =>
            state <= "1011010000";
            uut_rst <= '0';
          WHEN "1011010000" =>
            state <= "1011010001";
            uut_rst <= '0';
          WHEN "1011010001" =>
            state <= "1011010010";
            uut_rst <= '0';
          WHEN "1011010010" =>
            state <= "1011010011";
            uut_rst <= '0';
          WHEN "1011010011" =>
            state <= "1011010100";
            uut_rst <= '0';
          WHEN "1011010100" =>
            state <= "1011010101";
            uut_rst <= '0';
          WHEN "1011010101" =>
            state <= "1011010110";
            uut_rst <= '0';
          WHEN "1011010110" =>
            state <= "1011010111";
            uut_rst <= '0';
          WHEN "1011010111" =>
            state <= "1011011000";
            uut_rst <= '0';
          WHEN "1011011000" =>
            state <= "1011011001";
            uut_rst <= '0';
          WHEN "1011011001" =>
            state <= "1011011010";
            uut_rst <= '0';
          WHEN "1011011010" =>
            state <= "1011011011";
            uut_rst <= '0';
          WHEN "1011011011" =>
            state <= "1011011100";
            uut_rst <= '0';
          WHEN "1011011100" =>
            state <= "1011011101";
            uut_rst <= '0';
          WHEN "1011011101" =>
            state <= "1011011110";
            uut_rst <= '0';
          WHEN "1011011110" =>
            state <= "1011011111";
            uut_rst <= '0';
          WHEN "1011011111" =>
            state <= "1011100000";
            uut_rst <= '0';
          WHEN "1011100000" =>
            state <= "1011100001";
            uut_rst <= '0';
          WHEN "1011100001" =>
            state <= "1011100010";
            uut_rst <= '0';
          WHEN "1011100010" =>
            state <= "1011100011";
            uut_rst <= '0';
          WHEN "1011100011" =>
            state <= "1011100100";
            uut_rst <= '0';
          WHEN "1011100100" =>
            state <= "1011100101";
            uut_rst <= '0';
          WHEN "1011100101" =>
            state <= "1011100110";
            uut_rst <= '0';
          WHEN "1011100110" =>
            state <= "1011100111";
            uut_rst <= '0';
          WHEN "1011100111" =>
            state <= "1011101000";
            uut_rst <= '0';
          WHEN "1011101000" =>
            state <= "1011101001";
            uut_rst <= '0';
          WHEN "1011101001" =>
            state <= "1011101010";
            uut_rst <= '0';
          WHEN "1011101010" =>
            state <= "1011101011";
            uut_rst <= '0';
          WHEN "1011101011" =>
            state <= "1011101100";
            uut_rst <= '0';
          WHEN "1011101100" =>
            state <= "1011101101";
            uut_rst <= '0';
          WHEN "1011101101" =>
            state <= "1011101110";
            uut_rst <= '0';
          WHEN "1011101110" =>
            state <= "1011101111";
            uut_rst <= '0';
          WHEN "1011101111" =>
            state <= "1011110000";
            uut_rst <= '0';
          WHEN "1011110000" =>
            state <= "1011110001";
            uut_rst <= '0';
          WHEN "1011110001" =>
            state <= "1011110010";
            uut_rst <= '0';
          WHEN "1011110010" =>
            state <= "1011110011";
            uut_rst <= '0';
          WHEN "1011110011" =>
            state <= "1011110100";
            uut_rst <= '0';
          WHEN "1011110100" =>
            state <= "1011110101";
            uut_rst <= '0';
          WHEN "1011110101" =>
            state <= "1011110110";
            uut_rst <= '0';
          WHEN "1011110110" =>
            state <= "1011110111";
            uut_rst <= '0';
          WHEN "1011110111" =>
            state <= "1011111000";
            uut_rst <= '0';
          WHEN "1011111000" =>
            state <= "1011111001";
            uut_rst <= '0';
          WHEN "1011111001" =>
            state <= "1011111010";
            uut_rst <= '0';
          WHEN "1011111010" =>
            state <= "1011111011";
            uut_rst <= '0';
          WHEN "1011111011" =>
            state <= "1011111100";
            uut_rst <= '0';
          WHEN "1011111100" =>
            state <= "1011111101";
            uut_rst <= '0';
          WHEN "1011111101" =>
            state <= "1011111110";
            uut_rst <= '0';
          WHEN "1011111110" =>
            state <= "1011111111";
            uut_rst <= '0';
          WHEN "1011111111" =>
            state <= "1100000000";
            uut_rst <= '0';
          WHEN "1100000000" =>
            state <= "1100000001";
            uut_rst <= '0';
          WHEN "1100000001" =>
            state <= "1100000010";
            uut_rst <= '0';
          WHEN "1100000010" =>
            state <= "1100000011";
            uut_rst <= '0';
          WHEN "1100000011" =>
            state <= "1100000100";
            uut_rst <= '0';
          WHEN "1100000100" =>
            state <= "1100000101";
            uut_rst <= '0';
          WHEN "1100000101" =>
            state <= "1100000110";
            uut_rst <= '0';
          WHEN "1100000110" =>
            state <= "1100000111";
            uut_rst <= '0';
          WHEN "1100000111" =>
            state <= "1100001000";
            uut_rst <= '0';
          WHEN "1100001000" =>
            state <= "1100001001";
            uut_rst <= '0';
          WHEN "1100001001" =>
            state <= "1100001010";
            uut_rst <= '0';
          WHEN "1100001010" =>
            state <= "1100001011";
            uut_rst <= '0';
          WHEN "1100001011" =>
            state <= "1100001100";
            uut_rst <= '0';
          WHEN "1100001100" =>
            state <= "1100001101";
            uut_rst <= '0';
          WHEN "1100001101" =>
            state <= "1100001110";
            uut_rst <= '0';
          WHEN "1100001110" =>
            state <= "1100001111";
            uut_rst <= '0';
          WHEN "1100001111" =>
            state <= "1100010000";
            uut_rst <= '0';
          WHEN "1100010000" =>
            state <= "1100010001";
            uut_rst <= '0';
          WHEN "1100010001" =>
            state <= "1100010010";
            uut_rst <= '0';
          WHEN "1100010010" =>
            state <= "1100010011";
            uut_rst <= '0';
          WHEN "1100010011" =>
            state <= "1100010100";
            uut_rst <= '0';
          WHEN "1100010100" =>
            state <= "1100010101";
            uut_rst <= '0';
          WHEN "1100010101" =>
            state <= "1100010110";
            uut_rst <= '0';
          WHEN "1100010110" =>
            state <= "1100010111";
            uut_rst <= '0';
          WHEN "1100010111" =>
            state <= "1100011000";
            uut_rst <= '0';
          WHEN "1100011000" =>
            state <= "1100011001";
            uut_rst <= '0';
          WHEN "1100011001" =>
            state <= "1100011010";
            uut_rst <= '0';
          WHEN "1100011010" =>
            state <= "1100011011";
            uut_rst <= '0';
          WHEN "1100011011" =>
            state <= "1100011100";
            uut_rst <= '0';
          WHEN "1100011100" =>
            state <= "1100011101";
            uut_rst <= '0';
          WHEN "1100011101" =>
            state <= "1100011110";
            uut_rst <= '0';
          WHEN "1100011110" =>
            state <= "1100011111";
            uut_rst <= '0';
          WHEN "1100011111" =>
            state <= "1100100000";
            uut_rst <= '0';
          WHEN "1100100000" =>
            state <= "1100100001";
            uut_rst <= '0';
          WHEN "1100100001" =>
            state <= "1100100010";
            uut_rst <= '0';
          WHEN "1100100010" =>
            state <= "1100100011";
            uut_rst <= '0';
          WHEN "1100100011" =>
            state <= "1100100100";
            uut_rst <= '0';
          WHEN "1100100100" =>
            state <= "1100100101";
            uut_rst <= '0';
          WHEN "1100100101" =>
            state <= "1100100110";
            uut_rst <= '0';
          WHEN "1100100110" =>
            state <= "1100100111";
            uut_rst <= '0';
          WHEN "1100100111" =>
            state <= "1100101000";
            uut_rst <= '0';
          WHEN "1100101000" =>
            state <= "1100101001";
            uut_rst <= '0';
          WHEN "1100101001" =>
            state <= "1100101010";
            uut_rst <= '0';
          WHEN "1100101010" =>
            state <= "1100101011";
            uut_rst <= '0';
          WHEN "1100101011" =>
            state <= "1100101100";
            uut_rst <= '0';
          WHEN "1100101100" =>
            state <= "1100101101";
            uut_rst <= '0';
          WHEN "1100101101" =>
            state <= "1100101110";
            uut_rst <= '0';
          WHEN "1100101110" =>
            state <= "1100101111";
            uut_rst <= '0';
          WHEN "1100101111" =>
            state <= "1100110000";
            uut_rst <= '0';
          WHEN "1100110000" =>
            state <= "1100110001";
            uut_rst <= '0';
          WHEN "1100110001" =>
            state <= "1100110010";
            uut_rst <= '0';
          WHEN "1100110010" =>
            state <= "1100110011";
            uut_rst <= '0';
          WHEN "1100110011" =>
            state <= "1100110100";
            uut_rst <= '0';
          WHEN "1100110100" =>
            state <= "1100110101";
            uut_rst <= '0';
          WHEN "1100110101" =>
            state <= "1100110110";
            uut_rst <= '0';
          WHEN "1100110110" =>
            state <= "1100110111";
            uut_rst <= '0';
          WHEN "1100110111" =>
            state <= "1100111000";
            uut_rst <= '0';
          WHEN "1100111000" =>
            state <= "1100111001";
            uut_rst <= '0';
          WHEN "1100111001" =>
            state <= "1100111010";
            uut_rst <= '0';
          WHEN "1100111010" =>
            state <= "1100111011";
            uut_rst <= '0';
          WHEN "1100111011" =>
            state <= "1100111100";
            uut_rst <= '0';
          WHEN "1100111100" =>
            state <= "1100111101";
            uut_rst <= '0';
          WHEN "1100111101" =>
            state <= "1100111110";
            uut_rst <= '0';
          WHEN "1100111110" =>
            state <= "1100111111";
            uut_rst <= '0';
          WHEN "1100111111" =>
            state <= "1101000000";
            uut_rst <= '0';
          WHEN "1101000000" =>
            state <= "1101000001";
            uut_rst <= '0';
          WHEN "1101000001" =>
            state <= "1101000010";
            uut_rst <= '0';
          WHEN "1101000010" =>
            state <= "1101000011";
            uut_rst <= '0';
          WHEN "1101000011" =>
            state <= "1101000100";
            uut_rst <= '0';
          WHEN "1101000100" =>
            state <= "1101000101";
            uut_rst <= '0';
          WHEN "1101000101" =>
            state <= "1101000110";
            uut_rst <= '0';
          WHEN "1101000110" =>
            state <= "1101000111";
            uut_rst <= '0';
          WHEN "1101000111" =>
            state <= "1101001000";
            uut_rst <= '0';
          WHEN "1101001000" =>
            state <= "1101001001";
            uut_rst <= '0';
          WHEN "1101001001" =>
            state <= "1101001010";
            uut_rst <= '0';
          WHEN "1101001010" =>
            state <= "1101001011";
            uut_rst <= '0';
          WHEN "1101001011" =>
            state <= "1101001100";
            uut_rst <= '0';
          WHEN "1101001100" =>
            state <= "1101001101";
            uut_rst <= '0';
          WHEN "1101001101" =>
            state <= "1101001110";
            uut_rst <= '0';
          WHEN "1101001110" =>
            state <= "1101001111";
            uut_rst <= '0';
          WHEN "1101001111" =>
            state <= "1101010000";
            uut_rst <= '0';
          WHEN "1101010000" =>
            state <= "1101010001";
            uut_rst <= '0';
          WHEN OTHERS =>
            DONE <= '1';
            uut_rst <= '1';
        END CASE;
      END IF;
    END IF;
  END PROCESS;
END;
