/home/brandyn/fpga-image-registration/modules/./conv_3x3_derivatives/conv_3x3_derivatives.vhd