/home/brandyn/fpga-image-registration/modules/./vga_input_test/vga_timing_decode.vhd