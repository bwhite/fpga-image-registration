/home/brandyn/fpga-image-registration/modules/./fetch_stage/convert_2d_to_1d_coord.vhd