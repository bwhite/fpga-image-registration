/home/brandyn/fpga-image-registration/modules/./pyramid_stage/pyramid_stage.vhd