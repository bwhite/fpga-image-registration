/home/brandyn/fpga-image-registration/modules/./image_store_stage/memory_dump.vhd