/home/brandyn/fpga-image-registration/modules/./dvi_output_test/i2c_video_programmer.vhd