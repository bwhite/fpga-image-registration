/home/brandyn/fpga-image-registration/modules/./compute_stage/compute_stage.vhd