/home/brandyn/fpga-image-registration/modules/./dvi_output_test/dvi_video_test.vhd