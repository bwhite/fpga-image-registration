/home/brandyn/fpga-image-registration/modules/./zbt_ram_manager/zbt_controller.vhd