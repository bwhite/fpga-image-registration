/home/brandyn/fpga-image-registration/modules/./vga_input_test/vga_input.vhd