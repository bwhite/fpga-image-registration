/home/brandyn/fpga-image-registration/modules/./make_a_b_matrices/right_shifter.vhd