/home/brandyn/fpga-image-registration/modules/./fetch_stage/mem_addr_selector.vhd