LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
ENTITY compose_h_matrixT0_tb IS
PORT(
  CLK : IN STD_LOGIC;
  RST : IN STD_LOGIC;
  DONE : OUT STD_LOGIC;
  FAIL : OUT STD_LOGIC;
  FAIL_NUM : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END compose_h_matrixT0_tb;
ARCHITECTURE behavior OF compose_h_matrixT0_tb IS
  COMPONENT compose_h_matrix
  PORT(
    CLK : IN STD_LOGIC;
    RST : IN STD_LOGIC;
    VALID_IN : IN STD_LOGIC;
    H_0_0_I : IN STD_LOGIC_VECTOR(29 DOWNTO 0);
    H_1_0_I : IN STD_LOGIC_VECTOR(29 DOWNTO 0);
    H_0_1_I : IN STD_LOGIC_VECTOR(29 DOWNTO 0);
    H_1_1_I : IN STD_LOGIC_VECTOR(29 DOWNTO 0);
    H_0_2_I : IN STD_LOGIC_VECTOR(29 DOWNTO 0);
    H_1_2_I : IN STD_LOGIC_VECTOR(29 DOWNTO 0);
    P_0_0 : IN STD_LOGIC_VECTOR(29 DOWNTO 0);
    P_1_0 : IN STD_LOGIC_VECTOR(29 DOWNTO 0);
    P_0_1 : IN STD_LOGIC_VECTOR(29 DOWNTO 0);
    P_1_1 : IN STD_LOGIC_VECTOR(29 DOWNTO 0);
    P_0_2 : IN STD_LOGIC_VECTOR(29 DOWNTO 0);
    P_1_2 : IN STD_LOGIC_VECTOR(29 DOWNTO 0);
    VALID_OUT : OUT STD_LOGIC;
    H_0_0 : OUT STD_LOGIC_VECTOR(29 DOWNTO 0);
    H_1_0 : OUT STD_LOGIC_VECTOR(29 DOWNTO 0);
    H_0_1 : OUT STD_LOGIC_VECTOR(29 DOWNTO 0);
    H_1_1 : OUT STD_LOGIC_VECTOR(29 DOWNTO 0);
    H_0_2 : OUT STD_LOGIC_VECTOR(29 DOWNTO 0);
    H_1_2 : OUT STD_LOGIC_VECTOR(29 DOWNTO 0));
  END COMPONENT;
  SIGNAL uut_rst_wire, uut_rst : STD_LOGIC;
  SIGNAL state : STD_LOGIC_VECTOR(5 DOWNTO 0);
  -- UUT Input
  SIGNAL uut_valid_in : STD_LOGIC;
  SIGNAL uut_h_0_0_i, uut_h_1_0_i, uut_h_0_1_i, uut_h_1_1_i, uut_h_0_2_i, uut_h_1_2_i, uut_p_0_0, uut_p_1_0, uut_p_0_1, uut_p_1_1, uut_p_0_2, uut_p_1_2 : STD_LOGIC_VECTOR(29 DOWNTO 0);
  -- UUT Output
  SIGNAL uut_valid_out : STD_LOGIC;
  SIGNAL uut_h_0_0, uut_h_1_0, uut_h_0_1, uut_h_1_1, uut_h_0_2, uut_h_1_2 : STD_LOGIC_VECTOR(29 DOWNTO 0);
BEGIN
  uut_rst_wire <= RST OR uut_rst;
  uut :  compose_h_matrix PORT MAP (
    CLK => CLK,
    RST => uut_rst_wire,
    VALID_IN => uut_valid_in,
    H_0_0_I => uut_h_0_0_i,
    H_1_0_I => uut_h_1_0_i,
    H_0_1_I => uut_h_0_1_i,
    H_1_1_I => uut_h_1_1_i,
    H_0_2_I => uut_h_0_2_i,
    H_1_2_I => uut_h_1_2_i,
    P_0_0 => uut_p_0_0,
    P_1_0 => uut_p_1_0,
    P_0_1 => uut_p_0_1,
    P_1_1 => uut_p_1_1,
    P_0_2 => uut_p_0_2,
    P_1_2 => uut_p_1_2,
    VALID_OUT => uut_valid_out,
    H_0_0 => uut_h_0_0,
    H_1_0 => uut_h_1_0,
    H_0_1 => uut_h_0_1,
    H_1_1 => uut_h_1_1,
    H_0_2 => uut_h_0_2,
    H_1_2 => uut_h_1_2
  );
  PROCESS (CLK) IS
  BEGIN
    IF CLK'event AND CLK='1' THEN
      IF RST='1' THEN
        DONE <= '0';
        FAIL <= '0';
        uut_rst <= '1';
        FAIL_NUM <= (OTHERS => '0');
        state <= (OTHERS => '0');
      ELSE
        CASE state IS
          WHEN "000000" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000001010011111000001010001";
            uut_h_1_0_i <= "000000001110011011110100100111";
            uut_h_0_1_i <= "000000001110010101011101101110";
            uut_h_1_1_i <= "000000011011010000011010000110";
            uut_h_0_2_i <= "000000100100110000101011111000";
            uut_h_1_2_i <= "000000000011111010100000100000";
            uut_p_0_0 <= "000000010100001101000010010100";
            uut_p_1_0 <= "000000011000011110011011100011";
            uut_p_0_1 <= "000000011101011110011011000010";
            uut_p_1_1 <= "000000001100000001001101011011";
            uut_p_0_2 <= "000000001000011100111000101011";
            uut_p_1_2 <= "000000011100010011101101001011";
            state <= "000001";
            uut_rst <= '0';
          WHEN "000001" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000010100100111010101100001";
            uut_h_1_0_i <= "000000011110101010010010111000";
            uut_h_0_1_i <= "000000011011011011011011100001";
            uut_h_1_1_i <= "000000000000001011101101001011";
            uut_h_0_2_i <= "000000000101111110101111100011";
            uut_h_1_2_i <= "000000000110001111100110101000";
            uut_p_0_0 <= "000000001101011001111011011110";
            uut_p_1_0 <= "000000011001001101110010000011";
            uut_p_0_1 <= "000000000111100101100100100001";
            uut_p_1_1 <= "000000100011111001010010001100";
            uut_p_0_2 <= "000000010110001001001010001100";
            uut_p_1_2 <= "000000011000100010011011011101";
            state <= "000010";
            uut_rst <= '0';
          WHEN "000010" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000010101000001111101111110";
            uut_h_1_0_i <= "000000001000001000001101101110";
            uut_h_0_1_i <= "000000000000000010001100111001";
            uut_h_1_1_i <= "000000011100101011011000100001";
            uut_h_0_2_i <= "000000100110100110001111001010";
            uut_h_1_2_i <= "000000000101001011111000010011";
            uut_p_0_0 <= "000000100011101000001101011011";
            uut_p_1_0 <= "000000000101010101011101100000";
            uut_p_0_1 <= "000000100111110110010010110000";
            uut_p_1_1 <= "000000001101100101101110011101";
            uut_p_0_2 <= "000000011111100101001010101101";
            uut_p_1_2 <= "000000010110100110100010010101";
            state <= "000011";
            uut_rst <= '0';
          WHEN "000011" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000010101101101010110110011";
            uut_h_1_0_i <= "000000100011100110010100111010";
            uut_h_0_1_i <= "000000000001001000010111011000";
            uut_h_1_1_i <= "000000010110100101011011110001";
            uut_h_0_2_i <= "000000000100100000001100111110";
            uut_h_1_2_i <= "000000000001111000111001111101";
            uut_p_0_0 <= "000000001001011101111000010101";
            uut_p_1_0 <= "000000100011111111110111010110";
            uut_p_0_1 <= "000000100011111001101010000101";
            uut_p_1_1 <= "000000100111001001001010011000";
            uut_p_0_2 <= "000000011101101001110000110110";
            uut_p_1_2 <= "000000100110101001001101010100";
            state <= "000100";
            uut_rst <= '0';
          WHEN "000100" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000010010010101001101110111";
            uut_h_1_0_i <= "000000000100101110001101100110";
            uut_h_0_1_i <= "000000000001010000001001110011";
            uut_h_1_1_i <= "000000001001111001101010011110";
            uut_h_0_2_i <= "000000001010011100101000101110";
            uut_h_1_2_i <= "000000011101011101011000000011";
            uut_p_0_0 <= "000000001100100100001000101010";
            uut_p_1_0 <= "000000000111100101001101011011";
            uut_p_0_1 <= "000000011011011100101000110001";
            uut_p_1_1 <= "000000010100100001001101010000";
            uut_p_0_2 <= "000000010000001010000001011001";
            uut_p_1_2 <= "000000100101110100110111000110";
            state <= "000101";
            uut_rst <= '0';
          WHEN "000101" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000010001000001100110110111";
            uut_h_1_0_i <= "000000010001000001011011010000";
            uut_h_0_1_i <= "000000001111111101101001010001";
            uut_h_1_1_i <= "000000100010100011110011000101";
            uut_h_0_2_i <= "000000010111011100100100111110";
            uut_h_1_2_i <= "000000011101000101001111111110";
            uut_p_0_0 <= "000000000000100100111000110011";
            uut_p_1_0 <= "000000011110000111111001011000";
            uut_p_0_1 <= "000000001101010101010110011100";
            uut_p_1_1 <= "000000010010100011000001111010";
            uut_p_0_2 <= "000000001101010100101011101111";
            uut_p_1_2 <= "000000010010010000111011110101";
            state <= "000110";
            uut_rst <= '0';
          WHEN "000110" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000100110111000110111001011";
            uut_h_1_0_i <= "000000000001100110111011100011";
            uut_h_0_1_i <= "000000000100010111111010010001";
            uut_h_1_1_i <= "000000000100001100001001101111";
            uut_h_0_2_i <= "000000010010100101110101111011";
            uut_h_1_2_i <= "000000011010010011011101000100";
            uut_p_0_0 <= "000000010101000001011000001111";
            uut_p_1_0 <= "000000100111101010000010010011";
            uut_p_0_1 <= "000000001011010001111101000011";
            uut_p_1_1 <= "000000010111100101000001110010";
            uut_p_0_2 <= "000000010000010111010101110101";
            uut_p_1_2 <= "000000000000110110110001001011";
            state <= "000111";
            uut_rst <= '0';
          WHEN "000111" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000100110010010011101111010";
            uut_h_1_0_i <= "000000000101001011001000001001";
            uut_h_0_1_i <= "000000011001000111110011100111";
            uut_h_1_1_i <= "000000100010000010111000011111";
            uut_h_0_2_i <= "000000100001011111001011000110";
            uut_h_1_2_i <= "000000010000001100001111000011";
            uut_p_0_0 <= "000000100110001111000100100011";
            uut_p_1_0 <= "000000010000011001010100001101";
            uut_p_0_1 <= "000000011111010000101010110010";
            uut_p_1_1 <= "000000001010110111001011100100";
            uut_p_0_2 <= "000000100011101110001111010101";
            uut_p_1_2 <= "000000010101111000000010110110";
            state <= "001000";
            uut_rst <= '0';
          WHEN "001000" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000011001000111110010001110";
            uut_h_1_0_i <= "000000100000101001100100101010";
            uut_h_0_1_i <= "000000011111011101011110010110";
            uut_h_1_1_i <= "000000010010010010011111110001";
            uut_h_0_2_i <= "000000010110000100011011000000";
            uut_h_1_2_i <= "000000000111000110000111111000";
            uut_p_0_0 <= "000000000100110100011101101001";
            uut_p_1_0 <= "000000001101101111100101100100";
            uut_p_0_1 <= "000000010011010000011110111111";
            uut_p_1_1 <= "000000010110111111000101011001";
            uut_p_0_2 <= "000000001110010100011001110100";
            uut_p_1_2 <= "000000100000101000010000110001";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000100011001010110001110011100" OR uut_h_1_0 /= "000111011111010111111010010001" OR uut_h_0_1 /= "000011110000101010101110100101" OR uut_h_1_1 /= "000101111000100001111010111011" OR uut_h_0_2 /= "000100011011111101111100000011" OR uut_h_1_2 /= "000111000010101100100010001111" THEN
              FAIL <= '1';
              FAIL_NUM <= "000000";
              state <= "101001";
            ELSE
              state <= "001001";
            END IF;
            uut_rst <= '0';
          WHEN "001001" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000010100011101101110100100";
            uut_h_1_0_i <= "000000010011101000010110110111";
            uut_h_0_1_i <= "000000001101000001000011010000";
            uut_h_1_1_i <= "000000001010111111010000001101";
            uut_h_0_2_i <= "000000011000101011010011010111";
            uut_h_1_2_i <= "000000011010001001110100100111";
            uut_p_0_0 <= "000000000000111111010100010111";
            uut_p_1_0 <= "000000011100101101101000100100";
            uut_p_0_1 <= "000000001111111010011100011001";
            uut_p_1_1 <= "000000100000100001011010111100";
            uut_p_0_2 <= "000000100011000010001000011101";
            uut_p_1_2 <= "000000001100000000000101101110";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000111100011111110110101000111" OR uut_h_1_0 /= "000011001111110100000000010111" OR uut_h_0_1 /= "001000111010011110100100000110" OR uut_h_1_1 /= "000001110111100110000110000110" OR uut_h_0_2 /= "001000111010101111001011001110" OR uut_h_1_2 /= "000101011011111100111000010100" THEN
              FAIL <= '1';
              FAIL_NUM <= "000001";
              state <= "101001";
            ELSE
              state <= "001010";
            END IF;
            uut_rst <= '0';
          WHEN "001010" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000010100110011110110000111";
            uut_h_1_0_i <= "000000001100101011001101011101";
            uut_h_0_1_i <= "000000011111011111010001100111";
            uut_h_1_1_i <= "000000100010011000100001100011";
            uut_h_0_2_i <= "000000000000000001100001001000";
            uut_h_1_2_i <= "000000000100110001001010001000";
            uut_p_0_0 <= "000000000010000011011111111001";
            uut_p_1_0 <= "000000000100010010010001101111";
            uut_p_0_1 <= "000000000000101110001101100001";
            uut_p_1_1 <= "000000011101110100010111000001";
            uut_p_0_2 <= "000000010011001111111101001100";
            uut_p_1_2 <= "000000010100001101001101001111";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000101110110101111001000110011" OR uut_h_1_0 /= "000011011101010011010110101101" OR uut_h_0_1 /= "000110100011010000010000000000" OR uut_h_1_1 /= "000101100100110011110001100001" OR uut_h_0_2 /= "000101110011000100011100110101" OR uut_h_1_2 /= "000111001001101000000010100100" THEN
              FAIL <= '1';
              FAIL_NUM <= "000010";
              state <= "101001";
            ELSE
              state <= "001011";
            END IF;
            uut_rst <= '0';
          WHEN "001011" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000100101011100110010001110";
            uut_h_1_0_i <= "000000100001010000110010001101";
            uut_h_0_1_i <= "000000001011110000011100001001";
            uut_h_1_1_i <= "000000000101101011010101110001";
            uut_h_0_2_i <= "000000100111000110011110101000";
            uut_h_1_2_i <= "000000010001101011001011111011";
            uut_p_0_0 <= "000000000011001100001011101100";
            uut_p_1_0 <= "000000011100111111101111111011";
            uut_p_0_1 <= "000000010011010001100010010110";
            uut_p_1_1 <= "000000011101110000011111000111";
            uut_p_0_2 <= "000000000000111100001100100100";
            uut_p_1_2 <= "000000000100000011000111111001";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000001111011000110111011011111" OR uut_h_1_0 /= "001000111111000000100110011100" OR uut_h_0_1 /= "000110011011110011110111101000" OR uut_h_1_1 /= "010000111001000010011010001010" OR uut_h_0_2 /= "000101011100001101011010100111" OR uut_h_1_2 /= "001111000110000100100101011100" THEN
              FAIL <= '1';
              FAIL_NUM <= "000011";
              state <= "101001";
            ELSE
              state <= "001100";
            END IF;
            uut_rst <= '0';
          WHEN "001100" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000000110001110000000111000";
            uut_h_1_0_i <= "000000011000110000101110101001";
            uut_h_0_1_i <= "000000001010101100001100010011";
            uut_h_1_1_i <= "000000001100101100100111001001";
            uut_h_0_2_i <= "000000100010010001011001011111";
            uut_h_1_2_i <= "000000011011101101110011110111";
            uut_p_0_0 <= "000000010011110101111001101001";
            uut_p_1_0 <= "000000001010100111010001110001";
            uut_p_0_1 <= "000000100101010010010110100100";
            uut_p_1_1 <= "000000000000001101100100110001";
            uut_p_0_2 <= "000000010101100101001110110111";
            uut_p_1_2 <= "000000010001100100100000000111";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000001110111111010010101111010" OR uut_h_1_0 /= "000001000011001100100111101011" OR uut_h_0_1 /= "000100001000011011001110100011" OR uut_h_1_1 /= "000010100110011000100000011101" OR uut_h_0_2 /= "000010110110001110001010001001" OR uut_h_1_2 /= "000011111110110111001100110011" THEN
              FAIL <= '1';
              FAIL_NUM <= "000100";
              state <= "101001";
            ELSE
              state <= "001101";
            END IF;
            uut_rst <= '0';
          WHEN "001101" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000000111100000101101111010";
            uut_h_1_0_i <= "000000001000111100100000100100";
            uut_h_0_1_i <= "000000100000110010100101111100";
            uut_h_1_1_i <= "000000000110010100101100101110";
            uut_h_0_2_i <= "000000001111101011101011011101";
            uut_h_1_2_i <= "000000010100111001101101101000";
            uut_p_0_0 <= "000000011000110111100110010111";
            uut_p_1_0 <= "000000000101010110001010001010";
            uut_p_0_1 <= "000000010101100011110010110111";
            uut_p_1_1 <= "000000011011111011110101011010";
            uut_p_0_2 <= "000000010000111101100010101010";
            uut_p_1_2 <= "000000100010001110110111001011";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000011110101010101101101000101" OR uut_h_1_0 /= "001000001101011011010111111100" OR uut_h_0_1 /= "000100000101100010100101110101" OR uut_h_1_1 /= "000110110001111110011110001010" OR uut_h_0_2 /= "000100011010101001000011111110" OR uut_h_1_2 /= "000111001010000101010111011110" THEN
              FAIL <= '1';
              FAIL_NUM <= "000101";
              state <= "101001";
            ELSE
              state <= "001110";
            END IF;
            uut_rst <= '0';
          WHEN "001110" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000011111111111110001110001";
            uut_h_1_0_i <= "000000011100110100011001000101";
            uut_h_0_1_i <= "000000100000011000000011011001";
            uut_h_1_1_i <= "000000010111000111110111000010";
            uut_h_0_2_i <= "000000100010011100111101100101";
            uut_h_1_2_i <= "000000000111011100110001011011";
            uut_p_0_0 <= "000000010100110001101100111001";
            uut_p_1_0 <= "000000100101010100100000000100";
            uut_p_0_1 <= "000000011011010011010011011110";
            uut_p_1_1 <= "000000011011011010101011100000";
            uut_p_0_2 <= "000000001101110101101011101100";
            uut_p_1_2 <= "000000010111001100001111000101";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000111101111011110000010010001" OR uut_h_1_0 /= "000001100011111110111010000000" OR uut_h_0_1 /= "000100001110111001110010000100" OR uut_h_1_1 /= "000000111010011101110111111111" OR uut_h_0_2 /= "000101010010101010010110110000" OR uut_h_1_2 /= "000000101001010000011001110011" THEN
              FAIL <= '1';
              FAIL_NUM <= "000110";
              state <= "101001";
            ELSE
              state <= "001111";
            END IF;
            uut_rst <= '0';
          WHEN "001111" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000000101000010000000101100";
            uut_h_1_0_i <= "000000010010000000110010010100";
            uut_h_0_1_i <= "000000010010010100100001100010";
            uut_h_1_1_i <= "000000011101111110001001011100";
            uut_h_0_2_i <= "000000000110000000101110011001";
            uut_h_1_2_i <= "000000000101011000111011010011";
            uut_p_0_0 <= "000000000010001100110101101011";
            uut_p_1_0 <= "000000100111011000110010011001";
            uut_p_0_1 <= "000000001001110110001010000111";
            uut_p_1_1 <= "000000011001000101011101101101";
            uut_p_0_2 <= "000000000110100011001011111110";
            uut_p_1_2 <= "000000000101101011010010001000";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "001110101001111011110101111111" OR uut_h_1_0 /= "000101111010000000011001101100" OR uut_h_0_1 /= "001011011110111001100000010000" OR uut_h_1_1 /= "000100001001110001010100010111" OR uut_h_0_2 /= "001111100000001001100000110101" OR uut_h_1_2 /= "000111100000111110110111010010" THEN
              FAIL <= '1';
              FAIL_NUM <= "000111";
              state <= "101001";
            ELSE
              state <= "010000";
            END IF;
            uut_rst <= '0';
          WHEN "010000" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000011010000100111000101011";
            uut_h_1_0_i <= "000000000001010010111010101101";
            uut_h_0_1_i <= "000000010001011011111000011100";
            uut_h_1_1_i <= "000000011111001001001111101000";
            uut_h_0_2_i <= "000000011011010101001110101011";
            uut_h_1_2_i <= "000000001011110011010100101011";
            uut_p_0_0 <= "000000100100010110111100111011";
            uut_p_1_0 <= "000000100000100111000100100011";
            uut_p_0_1 <= "000000100001101111011011011100";
            uut_p_1_1 <= "000000011101000110110000001100";
            uut_p_0_2 <= "000000100110100101101000010010";
            uut_p_1_2 <= "000000100101001010010101111000";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000100010100101110101011111000" OR uut_h_1_0 /= "000011001100010110111110101101" OR uut_h_0_1 /= "001001011011011101100011100010" OR uut_h_1_1 /= "001000001100100100010111111110" OR uut_h_0_2 /= "001011001011001100000111010011" OR uut_h_1_2 /= "001000011011001110010101000100" THEN
              FAIL <= '1';
              FAIL_NUM <= "001000";
              state <= "101001";
            ELSE
              state <= "010001";
            END IF;
            uut_rst <= '0';
          WHEN "010001" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000001111011110000001000101";
            uut_h_1_0_i <= "000000011101001010011001000001";
            uut_h_0_1_i <= "000000100000111110001001111000";
            uut_h_1_1_i <= "000000000111100011100110011111";
            uut_h_0_2_i <= "000000010011011110000101110011";
            uut_h_1_2_i <= "000000000011010010100100100010";
            uut_p_0_0 <= "000000001000110100000110110100";
            uut_p_1_0 <= "000000011001011000011001001011";
            uut_p_0_1 <= "000000011001110011010001111100";
            uut_p_1_1 <= "000000000101000011101010010011";
            uut_p_0_2 <= "000000010111000110101101111100";
            uut_p_1_2 <= "000000010011011011100001100011";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000011000100111111100101110111" OR uut_h_1_0 /= "000010100111011101101111111110" OR uut_h_0_1 /= "000101110110011111010010011101" OR uut_h_1_1 /= "000101001110110111111111011000" OR uut_h_0_2 /= "000111001101010000001111001001" OR uut_h_1_2 /= "000110110011111101000000100110" THEN
              FAIL <= '1';
              FAIL_NUM <= "001001";
              state <= "101001";
            ELSE
              state <= "010010";
            END IF;
            uut_rst <= '0';
          WHEN "010010" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000100011011010101110110001";
            uut_h_1_0_i <= "000000001000100001111001111100";
            uut_h_0_1_i <= "000000100010010000010011101111";
            uut_h_1_1_i <= "000000010100100010101011000010";
            uut_h_0_2_i <= "000000010110011010101010111010";
            uut_h_1_2_i <= "000000001101101100101011011111";
            uut_p_0_0 <= "000000100011010111010000111010";
            uut_p_1_0 <= "000000011010000010010000110011";
            uut_p_0_1 <= "000000100111110011000011001000";
            uut_p_1_1 <= "000000100001010101100100001001";
            uut_p_0_2 <= "000000001010100110001010011111";
            uut_p_1_2 <= "000000100101001101000011111011";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000001011000110110100011100110" OR uut_h_1_0 /= "000001010110101100101001000100" OR uut_h_0_1 /= "000111011100111110101011111010" OR uut_h_1_1 /= "001000000101001100100111001101" OR uut_h_0_2 /= "001000000110011100110000011001" OR uut_h_1_2 /= "000111011010001001000100001011" THEN
              FAIL <= '1';
              FAIL_NUM <= "001010";
              state <= "101001";
            ELSE
              state <= "010011";
            END IF;
            uut_rst <= '0';
          WHEN "010011" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000000010011010100101010110";
            uut_h_1_0_i <= "000000000100110000110011101100";
            uut_h_0_1_i <= "000000010101011110001000101100";
            uut_h_1_1_i <= "000000001011010010010110110100";
            uut_h_0_2_i <= "000000010010100011111111010101";
            uut_h_1_2_i <= "000000000001111111010001100000";
            uut_p_0_0 <= "000000000111010011001011010000";
            uut_p_1_0 <= "000000001010100100100010011100";
            uut_p_0_1 <= "000000001000010101011100001011";
            uut_p_1_1 <= "000000100111011100111110000111";
            uut_p_0_2 <= "000000010100010011010110001010";
            uut_p_1_2 <= "000000011010100000001111101010";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000011100110001100001100011001" OR uut_h_1_0 /= "000010000111010111100000010101" OR uut_h_0_1 /= "001000010111110101001110010010" OR uut_h_1_1 /= "000110010101000001001010110101" OR uut_h_0_2 /= "000001010000100000111000101101" OR uut_h_1_2 /= "000000101100110011110111010100" THEN
              FAIL <= '1';
              FAIL_NUM <= "001011";
              state <= "101001";
            ELSE
              state <= "010100";
            END IF;
            uut_rst <= '0';
          WHEN "010100" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000001011101111011000011111";
            uut_h_1_0_i <= "000000010110010011000010101101";
            uut_h_0_1_i <= "000000000111010110111110001011";
            uut_h_1_1_i <= "000000000111010110100110001101";
            uut_h_0_2_i <= "000000100001011100110111111111";
            uut_h_1_2_i <= "000000010000101000111001101100";
            uut_p_0_0 <= "000000011100011010100010111101";
            uut_p_1_0 <= "000000011001110101010001100000";
            uut_p_0_1 <= "000000001010111010101110111110";
            uut_p_1_1 <= "000000001100000100001101010110";
            uut_p_0_2 <= "000000000101010100000101010110";
            uut_p_1_2 <= "000000100100100101101000100010";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000001110110011011101001000110" OR uut_h_1_0 /= "000100111001000010101010011011" OR uut_h_0_1 /= "000001110101000100111000001110" OR uut_h_1_1 /= "000111001110111110111000000111" OR uut_h_0_2 /= "000011000011010011000011101111" OR uut_h_1_2 /= "000110010110011101010110100101" THEN
              FAIL <= '1';
              FAIL_NUM <= "001100";
              state <= "101001";
            ELSE
              state <= "010101";
            END IF;
            uut_rst <= '0';
          WHEN "010101" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000000001010001010001011100";
            uut_h_1_0_i <= "000000001110111111110011101011";
            uut_h_0_1_i <= "000000100010001011110011100110";
            uut_h_1_1_i <= "000000011011011100100010110011";
            uut_h_0_2_i <= "000000010001100111110010101000";
            uut_h_1_2_i <= "000000000011000111010111011111";
            uut_p_0_0 <= "000000011010000001111000010111";
            uut_p_1_0 <= "000000010011011110100100000010";
            uut_p_0_1 <= "000000001001011100101101101101";
            uut_p_1_1 <= "000000011000011101101101101000";
            uut_p_0_2 <= "000000011000100110001110100111";
            uut_p_1_2 <= "000000011101000110010111101110";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000010110101000011001100100010" OR uut_h_1_0 /= "000010000000001000100101111010" OR uut_h_0_1 /= "001000011010111101111101110100" OR uut_h_1_1 /= "000010111000110000000011011100" OR uut_h_0_2 /= "001010000000101000010010011000" OR uut_h_1_2 /= "000011001100111111111010001100" THEN
              FAIL <= '1';
              FAIL_NUM <= "001101";
              state <= "101001";
            ELSE
              state <= "010110";
            END IF;
            uut_rst <= '0';
          WHEN "010110" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000100111100010011110011101";
            uut_h_1_0_i <= "000000011110011100011110100100";
            uut_h_0_1_i <= "000000100010010111011100110101";
            uut_h_1_1_i <= "000000011000111101111010011101";
            uut_h_0_2_i <= "000000010010111011010001100100";
            uut_h_1_2_i <= "000000010001111100011010101010";
            uut_p_0_0 <= "000000011111011001101101100111";
            uut_p_1_0 <= "000000100010000010001111001011";
            uut_p_0_1 <= "000000011010110110101011101101";
            uut_p_1_1 <= "000000001101110110100101101111";
            uut_p_0_2 <= "000000000111100100000110010001";
            uut_p_1_2 <= "000000001100101011101101000010";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "001110101000100001110000101010" OR uut_h_1_0 /= "001011011010110110100000100101" OR uut_h_0_1 /= "001101110000100110011011110100" OR uut_h_1_1 /= "001011000110011000000000110100" OR uut_h_0_2 /= "001001110111010001000001011110" OR uut_h_1_2 /= "000111011010111110101100101001" THEN
              FAIL <= '1';
              FAIL_NUM <= "001110";
              state <= "101001";
            ELSE
              state <= "010111";
            END IF;
            uut_rst <= '0';
          WHEN "010111" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000010011001011000111000101";
            uut_h_1_0_i <= "000000010001111011010111100001";
            uut_h_0_1_i <= "000000100010010011011011010111";
            uut_h_1_1_i <= "000000011010010100110101010101";
            uut_h_0_2_i <= "000000011110001000010100000101";
            uut_h_1_2_i <= "000000100000100010101000000101";
            uut_p_0_0 <= "000000011000101100100001100110";
            uut_p_1_0 <= "000000000110001110100001001001";
            uut_p_0_1 <= "000000001100100110000010001101";
            uut_p_1_1 <= "000000011011100110110100110010";
            uut_p_0_2 <= "000000011011000011101001001000";
            uut_p_1_2 <= "000000001010000001001001011001";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000101101110010101100101100000" OR uut_h_1_0 /= "001001100010000011101111010100" OR uut_h_0_1 /= "000011111110100011111001010110" OR uut_h_1_1 /= "000111010000100110000001001000" OR uut_h_0_2 /= "000001001010011111000100110111" OR uut_h_1_2 /= "000010010101011100001011001010" THEN
              FAIL <= '1';
              FAIL_NUM <= "001111";
              state <= "101001";
            ELSE
              state <= "011000";
            END IF;
            uut_rst <= '0';
          WHEN "011000" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000000001110010010001001001";
            uut_h_1_0_i <= "000000100111011000001010001011";
            uut_h_0_1_i <= "000000100000000111010110110101";
            uut_h_1_1_i <= "000000011101110101111101100000";
            uut_h_0_2_i <= "000000010000101100011000111010";
            uut_h_1_2_i <= "000000010000010000000111001101";
            uut_p_0_0 <= "000000010100111101010011100111";
            uut_p_1_0 <= "000000001111001000001001011010";
            uut_p_0_1 <= "000000001111010010111111111100";
            uut_p_1_1 <= "000000011001000010011011101111";
            uut_p_0_2 <= "000000011011110100000001101001";
            uut_p_1_2 <= "000000011000110110010010010101";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "001011110110010101111010011110" OR uut_h_1_0 /= "001000010011010111101101010001" OR uut_h_0_1 /= "001010110101101010001001101101" OR uut_h_1_1 /= "000111011011000110000011100110" OR uut_h_0_2 /= "001101010110011010101001001101" OR uut_h_1_2 /= "001001100111011111001100000001" THEN
              FAIL <= '1';
              FAIL_NUM <= "010000";
              state <= "101001";
            ELSE
              state <= "011001";
            END IF;
            uut_rst <= '0';
          WHEN "011001" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000010011101110000000111110";
            uut_h_1_0_i <= "000000001111011001011110010111";
            uut_h_0_1_i <= "000000100000000101001000100001";
            uut_h_1_1_i <= "000000010011110101001011110100";
            uut_h_0_2_i <= "000000100010011011100010111101";
            uut_h_1_2_i <= "000000010101010010011110110110";
            uut_p_0_0 <= "000000100110010100000100011110";
            uut_p_1_0 <= "000000100100010110010011011010";
            uut_p_0_1 <= "000000000000001011110111010000";
            uut_p_1_1 <= "000000001111010000111101100100";
            uut_p_0_2 <= "000000011100111101001000001100";
            uut_p_1_2 <= "000000010010101001000010000110";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000111100110100110001001101100" OR uut_h_1_0 /= "000011100000011010100000111010" OR uut_h_0_1 /= "000100011010111011100100110110" OR uut_h_1_1 /= "000110001011010100011100100111" OR uut_h_0_2 /= "001000000110011111011101011110" OR uut_h_1_2 /= "000110011101100110001110001010" THEN
              FAIL <= '1';
              FAIL_NUM <= "010001";
              state <= "101001";
            ELSE
              state <= "011010";
            END IF;
            uut_rst <= '0';
          WHEN "011010" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000000111000011110110000110";
            uut_h_1_0_i <= "000000011110010111000111100100";
            uut_h_0_1_i <= "000000001110110101111111000111";
            uut_h_1_1_i <= "000000100001100111010001111011";
            uut_h_0_2_i <= "000000011010101110011111110100";
            uut_h_1_2_i <= "000000011110100011000111110100";
            uut_p_0_0 <= "000000011010111010001011010010";
            uut_p_1_0 <= "000000010011011001001111010011";
            uut_p_0_1 <= "000000001000000011000101110101";
            uut_p_1_1 <= "000000010010010010010000110000";
            uut_p_0_2 <= "000000100010011011011101010001";
            uut_p_1_2 <= "000000000011111100001001000110";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "010000110000001010100001101110" OR uut_h_1_0 /= "000110100010001110100010100000" OR uut_h_0_1 /= "010011111011101111101100101111" OR uut_h_1_1 /= "001000000000001000011100111101" OR uut_h_0_2 /= "001101001111010001100100100010" OR uut_h_1_2 /= "000110111001000000100011110011" THEN
              FAIL <= '1';
              FAIL_NUM <= "010010";
              state <= "101001";
            ELSE
              state <= "011011";
            END IF;
            uut_rst <= '0';
          WHEN "011011" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000000010010000001010100101";
            uut_h_1_0_i <= "000000100101011001011111101010";
            uut_h_0_1_i <= "000000100111100000111110011001";
            uut_h_1_1_i <= "000000100010011001100011111110";
            uut_h_0_2_i <= "000000001110011101000000010111";
            uut_h_1_2_i <= "000000000110110011011111110111";
            uut_p_0_0 <= "000000100010011010001001100000";
            uut_p_1_0 <= "000000001101001111100001010111";
            uut_p_0_1 <= "000000000010111101100100100100";
            uut_p_1_1 <= "000000000100100110000010111100";
            uut_p_0_2 <= "000000001110010000111000111100";
            uut_p_1_2 <= "000000011101101111010000000100";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000001111010010011001000011010" OR uut_h_1_0 /= "000001001101000010011110001011" OR uut_h_0_1 /= "000110110001100110111000100101" OR uut_h_1_1 /= "000011110010011111101110101001" OR uut_h_0_2 /= "000101000111100111000111001111" OR uut_h_1_2 /= "000011000111111010000001011010" THEN
              FAIL <= '1';
              FAIL_NUM <= "010011";
              state <= "101001";
            ELSE
              state <= "011100";
            END IF;
            uut_rst <= '0';
          WHEN "011100" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000001010100100110100100100";
            uut_h_1_0_i <= "000000001001011100101100010000";
            uut_h_0_1_i <= "000000100101100000100100110101";
            uut_h_1_1_i <= "000000001011111111010101100111";
            uut_h_0_2_i <= "000000000110100100111001101000";
            uut_h_1_2_i <= "000000011110001110110010011111";
            uut_p_0_0 <= "000000000011101110110010001010";
            uut_p_1_0 <= "000000011011010000000011110101";
            uut_p_0_1 <= "000000001001110010001001101101";
            uut_p_1_1 <= "000000010000001000110110010101";
            uut_p_0_2 <= "000000100110000111111010110101";
            uut_p_1_2 <= "000000000101011110101110111100";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000100000101110110010110001101" OR uut_h_1_0 /= "000110011011110000110111110000" OR uut_h_0_1 /= "000001101100011111000000010010" OR uut_h_1_1 /= "000010100110000101000100110110" OR uut_h_0_2 /= "000011000111010001001011100100" OR uut_h_1_2 /= "000011010010011001100001001001" THEN
              FAIL <= '1';
              FAIL_NUM <= "010100";
              state <= "101001";
            ELSE
              state <= "011101";
            END IF;
            uut_rst <= '0';
          WHEN "011101" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000100100110100000110000101";
            uut_h_1_0_i <= "000000011110000111011001010011";
            uut_h_0_1_i <= "000000100101000110111011111101";
            uut_h_1_1_i <= "000000000111011010101011111110";
            uut_h_0_2_i <= "000000011001001100001011000111";
            uut_h_1_2_i <= "000000000111111111000111100000";
            uut_p_0_0 <= "000000100000110110111010010010";
            uut_p_1_0 <= "000000001100001110100110111011";
            uut_p_0_1 <= "000000000000011001011100001001";
            uut_p_1_1 <= "000000011000101010001100111100";
            uut_p_0_2 <= "000000100100111100111011100000";
            uut_p_1_2 <= "000000100101000000111101010000";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000101011101011100010010001011" OR uut_h_1_0 /= "000111001110011110001011011010" OR uut_h_0_1 /= "000110101000001001011111011100" OR uut_h_1_1 /= "000110010110100100101110000101" OR uut_h_0_2 /= "001000010010100111011010001111" OR uut_h_1_2 /= "001001001010111001000001000110" THEN
              FAIL <= '1';
              FAIL_NUM <= "010101";
              state <= "101001";
            ELSE
              state <= "011110";
            END IF;
            uut_rst <= '0';
          WHEN "011110" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000011000100110110011000110";
            uut_h_1_0_i <= "000000011000111111011010111110";
            uut_h_0_1_i <= "000000001011011110100001110011";
            uut_h_1_1_i <= "000000011010001010100001001100";
            uut_h_0_2_i <= "000000001001110001100001000000";
            uut_h_1_2_i <= "000000000100100110101100011111";
            uut_p_0_0 <= "000000100101000100000011110010";
            uut_p_1_0 <= "000000010001111000110110010011";
            uut_p_0_1 <= "000000011111000001010110001101";
            uut_p_1_1 <= "000000010100110111101111000111";
            uut_p_0_2 <= "000000001111111000100010100111";
            uut_p_1_2 <= "000000011100100100010110000110";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "010010110101100111110010110110" OR uut_h_1_0 /= "001110000110111001010000111111" OR uut_h_0_1 /= "001100000000111011101011101010" OR uut_h_1_1 /= "001001000101101110100010001000" OR uut_h_0_2 /= "000110000010011001001111100000" OR uut_h_1_2 /= "000100100011011010101001100110" THEN
              FAIL <= '1';
              FAIL_NUM <= "010110";
              state <= "101001";
            ELSE
              state <= "011111";
            END IF;
            uut_rst <= '0';
          WHEN "011111" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000010011001110000011000110";
            uut_h_1_0_i <= "000000010100110111110101001001";
            uut_h_0_1_i <= "000000011000010111011101011111";
            uut_h_1_1_i <= "000000000011001011010111010011";
            uut_h_0_2_i <= "000000011100010101110110010001";
            uut_h_1_2_i <= "000000000001011101000110111001";
            uut_p_0_0 <= "000000011111000111100000100010";
            uut_p_1_0 <= "000000000110110110011101011000";
            uut_p_0_1 <= "000000011011111001000010111011";
            uut_p_1_1 <= "000000000101011001111101101101";
            uut_p_0_2 <= "000000001001111100010000001100";
            uut_p_1_2 <= "000000010110010011101110111101";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000101010111100011011101111010" OR uut_h_1_0 /= "000100101111010101000111011011" OR uut_h_0_1 /= "001001010010001111011110011101" OR uut_h_1_1 /= "000111011100010001011011010100" OR uut_h_0_2 /= "000111001101010110000010000111" OR uut_h_1_2 /= "000110010110111011111111111000" THEN
              FAIL <= '1';
              FAIL_NUM <= "010111";
              state <= "101001";
            ELSE
              state <= "100000";
            END IF;
            uut_rst <= '0';
          WHEN "100000" =>
            uut_valid_in <= '1';
            uut_h_0_0_i <= "000000000100111111101110101011";
            uut_h_1_0_i <= "000000000000111001101011011001";
            uut_h_0_1_i <= "000000010000100010100101011001";
            uut_h_1_1_i <= "000000000100101011100000111100";
            uut_h_0_2_i <= "000000010011100000011111100000";
            uut_h_1_2_i <= "000000010010000000001110011000";
            uut_p_0_0 <= "000000011010110000010001000011";
            uut_p_1_0 <= "000000011010110110001111001111";
            uut_p_0_1 <= "000000001010111010100000001110";
            uut_p_1_1 <= "000000011001001111000000010001";
            uut_p_0_2 <= "000000100111101110011111100100";
            uut_p_1_2 <= "000000100010011100011000000111";
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000100000101100111011001110000" OR uut_h_1_0 /= "001001111110010110111010000101" OR uut_h_0_1 /= "000110011111101101000000000101" OR uut_h_1_1 /= "001010100010110010000101000111" OR uut_h_0_2 /= "000110111000100001011011100101" OR uut_h_1_2 /= "001110100110101000001001011000" THEN
              FAIL <= '1';
              FAIL_NUM <= "011000";
              state <= "101001";
            ELSE
              state <= "100001";
            END IF;
            uut_rst <= '0';
          WHEN "100001" =>
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "001111000000110010010011101000" OR uut_h_1_0 /= "001010001111011001000000000010" OR uut_h_0_1 /= "000011110110101011100010001101" OR uut_h_1_1 /= "000010011000110010011001111101" OR uut_h_0_2 /= "001001101010111010110100001000" OR uut_h_1_2 /= "000110101101000011010001001110" THEN
              FAIL <= '1';
              FAIL_NUM <= "011001";
              state <= "101001";
            ELSE
              state <= "100010";
            END IF;
            uut_rst <= '0';
          WHEN "100010" =>
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000011101110111011100010011100" OR uut_h_1_0 /= "001011011110011101000010010101" OR uut_h_0_1 /= "000010100100000111101100111000" OR uut_h_1_1 /= "000110101101011111110101101110" OR uut_h_0_2 /= "000010110001100000001000010111" OR uut_h_1_2 /= "001001101011011010101010110110" THEN
              FAIL <= '1';
              FAIL_NUM <= "011010";
              state <= "101001";
            ELSE
              state <= "100011";
            END IF;
            uut_rst <= '0';
          WHEN "100011" =>
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000100101100011001010000100111" OR uut_h_1_0 /= "001101100111001011011110100000" OR uut_h_0_1 /= "000001011110000111001010001000" OR uut_h_1_1 /= "000010000110011010010101000011" OR uut_h_0_2 /= "001001101010000100111000110001" OR uut_h_1_2 /= "001100010001000001001000100111" THEN
              FAIL <= '1';
              FAIL_NUM <= "011011";
              state <= "101001";
            ELSE
              state <= "100100";
            END IF;
            uut_rst <= '0';
          WHEN "100100" =>
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "001000010010110011100100100000" OR uut_h_1_0 /= "000010110100111111011000100110" OR uut_h_0_1 /= "000101100010011001011100001011" OR uut_h_1_1 /= "000010001110111101110010001001" OR uut_h_0_2 /= "000100110110111100001101001111" OR uut_h_1_2 /= "000011110011001011111011000010" THEN
              FAIL <= '1';
              FAIL_NUM <= "011100";
              state <= "101001";
            ELSE
              state <= "100101";
            END IF;
            uut_rst <= '0';
          WHEN "100101" =>
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "001100111111101100111011000010" OR uut_h_1_0 /= "001000011100000111011100111101" OR uut_h_0_1 /= "000111010000110110100010010011" OR uut_h_1_1 /= "000001100001011011110100001100" OR uut_h_0_2 /= "010101110000001001100000001001" OR uut_h_1_2 /= "001010111101101010111101001100" THEN
              FAIL <= '1';
              FAIL_NUM <= "011101";
              state <= "101001";
            ELSE
              state <= "100110";
            END IF;
            uut_rst <= '0';
          WHEN "100110" =>
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "001000101110101001011010111111" OR uut_h_1_0 /= "001010111001001001000111111011" OR uut_h_0_1 /= "000111110101011011000100010101" OR uut_h_1_1 /= "001010010100101010001100100101" OR uut_h_0_2 /= "000101110001001000000101110011" OR uut_h_1_2 /= "001001000000110011100101111111" THEN
              FAIL <= '1';
              FAIL_NUM <= "011110";
              state <= "101001";
            ELSE
              state <= "100111";
            END IF;
            uut_rst <= '0';
          WHEN "100111" =>
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000101111110011111110001100000" OR uut_h_1_0 /= "000101001111101000010101111101" OR uut_h_0_1 /= "000101001101111000110100111011" OR uut_h_1_1 /= "000100101011101010101101010111" OR uut_h_0_2 /= "000110001011101010100100011011" OR uut_h_1_2 /= "000010001100101001100000101011" THEN
              FAIL <= '1';
              FAIL_NUM <= "011111";
              state <= "101001";
            ELSE
              state <= "101000";
            END IF;
            uut_rst <= '0';
          WHEN "101000" =>
            IF uut_valid_out /= '1' OR uut_h_0_0 /= "000100100000110111001100101001" OR uut_h_1_0 /= "000001001010111000001010101111" OR uut_h_0_1 /= "000011101011111101001010111100" OR uut_h_1_1 /= "000000111111111101110010110100" OR uut_h_0_2 /= "000110010011100101111101011010" OR uut_h_1_2 /= "000001110100100000000010110110" THEN
              FAIL <= '1';
              FAIL_NUM <= "100000";
              state <= "101001";
            ELSE
              state <= "101001";
            END IF;
            uut_rst <= '0';
          WHEN OTHERS =>
            DONE <= '1';
            uut_rst <= '1';
        END CASE;
      END IF;
    END IF;
  END PROCESS;
END;
