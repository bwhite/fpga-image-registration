/home/brandyn/fpga-image-registration/modules/./smooth_stage/pixel_conv_buf_3x3.vhd