/home/brandyn/fpga-image-registration/modules/./sum_a_b_matrices/sum_a_b_matrices.vhd