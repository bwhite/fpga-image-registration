/home/brandyn/fpga-image-registration/modules/./dvi_output_test/vga_timing_generator.vhd