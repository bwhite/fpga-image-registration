/home/brandyn/fpga-image-registration/modules/./dvi_output_test/const_test.vhd