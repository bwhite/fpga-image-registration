/home/brandyn/fpga-image-registration/modules/./unscale_h_matrix/unscale_h_matrix.vhd