/home/brandyn/fpga-image-registration/modules/./image_store_stage/image_store_display_test.vhd