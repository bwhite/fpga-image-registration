/home/brandyn/fpga-image-registration/modules/./image_store_stage/pixel_memory_controller.vhd