/home/brandyn/fpga-image-registration/modules/./affine_coord_transform/affine_coord_transform.vhd