/home/brandyn/fpga-image-registration/modules/./fetch_stage/img1_compute_mem_addr.vhd