../pixel_memory_test/pixel_memory_controller.vhd