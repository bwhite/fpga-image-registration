/home/brandyn/fpga-image-registration/modules/./conv_pixel_ordering/conv_pixel_ordering.vhd