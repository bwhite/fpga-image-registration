library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity make_h_matrix is
    Port ( CLK : in  STD_LOGIC;
           RST : in  STD_LOGIC);
end make_h_matrix;

architecture Behavioral of make_h_matrix is

begin


end Behavioral;

