LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
ENTITY unscale_h_matrixT0_tb IS
PORT(
  CLK : IN STD_LOGIC;
  RST : IN STD_LOGIC;
  DONE : OUT STD_LOGIC;
  FAIL : OUT STD_LOGIC;
  FAIL_NUM : OUT STD_LOGIC_VECTOR(5 DOWNTO 0));
END unscale_h_matrixT0_tb;
ARCHITECTURE behavior OF unscale_h_matrixT0_tb IS
  COMPONENT unscale_h_matrix
  PORT(
    CLK : IN STD_LOGIC;
    RST : IN STD_LOGIC;
    H_0_0_I : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    H_0_1_I : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    H_0_2_I : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    H_1_0_I : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    H_1_1_I : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    H_1_2_I : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    COORD_TRANS : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    INPUT_VALID : IN STD_LOGIC;
    H_0_0 : OUT STD_LOGIC_VECTOR(29 DOWNTO 0);
    H_0_1 : OUT STD_LOGIC_VECTOR(29 DOWNTO 0);
    H_0_2 : OUT STD_LOGIC_VECTOR(29 DOWNTO 0);
    H_1_0 : OUT STD_LOGIC_VECTOR(29 DOWNTO 0);
    H_1_1 : OUT STD_LOGIC_VECTOR(29 DOWNTO 0);
    H_1_2 : OUT STD_LOGIC_VECTOR(29 DOWNTO 0);
    OUTPUT_VALID : OUT STD_LOGIC);
  END COMPONENT;
  SIGNAL uut_rst_wire, uut_rst : STD_LOGIC;
  SIGNAL state : STD_LOGIC_VECTOR(5 DOWNTO 0);
  -- UUT Input
  SIGNAL uut_input_valid : STD_LOGIC;
  SIGNAL uut_h_0_0_i, uut_h_0_1_i, uut_h_0_2_i, uut_h_1_0_i, uut_h_1_1_i, uut_h_1_2_i : STD_LOGIC_VECTOR(26 DOWNTO 0);
  SIGNAL uut_coord_trans : STD_LOGIC_VECTOR(11 DOWNTO 0);
  -- UUT Output
  SIGNAL uut_output_valid : STD_LOGIC;
  SIGNAL uut_h_0_0, uut_h_0_1, uut_h_0_2, uut_h_1_0, uut_h_1_1, uut_h_1_2 : STD_LOGIC_VECTOR(29 DOWNTO 0);
BEGIN
  uut_rst_wire <= RST OR uut_rst;
  uut :  unscale_h_matrix PORT MAP (
    CLK => CLK,
    RST => uut_rst_wire,
    H_0_0_I => uut_h_0_0_i,
    H_0_1_I => uut_h_0_1_i,
    H_0_2_I => uut_h_0_2_i,
    H_1_0_I => uut_h_1_0_i,
    H_1_1_I => uut_h_1_1_i,
    H_1_2_I => uut_h_1_2_i,
    COORD_TRANS => uut_coord_trans,
    INPUT_VALID => uut_input_valid,
    H_0_0 => uut_h_0_0,
    H_0_1 => uut_h_0_1,
    H_0_2 => uut_h_0_2,
    H_1_0 => uut_h_1_0,
    H_1_1 => uut_h_1_1,
    H_1_2 => uut_h_1_2,
    OUTPUT_VALID => uut_output_valid
  );
  PROCESS (CLK) IS
  BEGIN
    IF CLK'event AND CLK='1' THEN
      IF RST='1' THEN
        DONE <= '0';
        FAIL <= '0';
        uut_rst <= '1';
        FAIL_NUM <= (OTHERS => '0');
        state <= (OTHERS => '0');
      ELSE
        CASE state IS
          WHEN "000000" =>
            uut_h_0_0_i <= "000000000000010111101110000";
            uut_h_0_1_i <= "111111110010111101001110100";
            uut_h_0_2_i <= "111111110011000101110100110";
            uut_h_1_0_i <= "000000000010000000000011100";
            uut_h_1_1_i <= "000000001011111011000010101";
            uut_h_1_2_i <= "000000001011000100010111100";
            uut_coord_trans <= "111110011110";
            uut_input_valid <= '1';
            state <= "000001";
            uut_rst <= '0';
          WHEN "000001" =>
            uut_h_0_0_i <= "000000000000110000100000001";
            uut_h_0_1_i <= "000000000100110001110001010";
            uut_h_0_2_i <= "000000000100001110001010111";
            uut_h_1_0_i <= "000000000100110011111010000";
            uut_h_1_1_i <= "000000001000011010010100101";
            uut_h_1_2_i <= "111111111000111001110000110";
            uut_coord_trans <= "111111110001";
            uut_input_valid <= '1';
            state <= "000010";
            uut_rst <= '0';
          WHEN "000010" =>
            uut_h_0_0_i <= "000000000100001101100100000";
            uut_h_0_1_i <= "111111111100110100110101110";
            uut_h_0_2_i <= "111111110010111001000110110";
            uut_h_1_0_i <= "000000001010101010111100001";
            uut_h_1_1_i <= "000000000001101111000111010";
            uut_h_1_2_i <= "000000000111110100011111100";
            uut_coord_trans <= "111111110001";
            uut_input_valid <= '1';
            state <= "000011";
            uut_rst <= '0';
          WHEN "000011" =>
            uut_h_0_0_i <= "111111110001001100010100000";
            uut_h_0_1_i <= "000000001101000110111011000";
            uut_h_0_2_i <= "111111111000001010010001101";
            uut_h_1_0_i <= "000000001111001110011011110";
            uut_h_1_1_i <= "111111111100010000111001000";
            uut_h_1_2_i <= "000000001101000101101110111";
            uut_coord_trans <= "111111101011";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000000010111101110000" OR uut_h_0_1 /= "111111111110010111101001110100" OR uut_h_0_2 /= "111101001110110001000001001010" OR uut_h_1_0 /= "000000000000010000000000011100" OR uut_h_1_1 /= "000000000001011111011000010101" OR uut_h_1_2 /= "111111110100101010100000011101" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "000000";
              state <= "111110";
            ELSE
              state <= "000100";
            END IF;
            uut_rst <= '0';
          WHEN "000100" =>
            uut_h_0_0_i <= "000000000100000000000010100";
            uut_h_0_1_i <= "111111110110110110100111001";
            uut_h_0_2_i <= "111111110111100001100001110";
            uut_h_1_0_i <= "000000000010001010011100000";
            uut_h_1_1_i <= "111111110000000111111001110";
            uut_h_1_2_i <= "111111110111110101011110111";
            uut_coord_trans <= "111111011000";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000000110000100000001" OR uut_h_0_1 /= "000000000000100110001110001010" OR uut_h_0_2 /= "111111110110101101111001101010" OR uut_h_1_0 /= "000000000000100110011111010000" OR uut_h_1_1 /= "000000000001000011010010100101" OR uut_h_1_2 /= "111111111100100000100011110100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "000001";
              state <= "111110";
            ELSE
              state <= "000101";
            END IF;
            uut_rst <= '0';
          WHEN "000101" =>
            uut_h_0_0_i <= "000000001010011010110111110";
            uut_h_0_1_i <= "111111111100100000010110010";
            uut_h_0_2_i <= "000000000100000000010101101";
            uut_h_1_0_i <= "000000001100010001110010110";
            uut_h_1_1_i <= "000000001001101001000110100";
            uut_h_1_2_i <= "000000000110010111100001011";
            uut_coord_trans <= "000000000110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000100001101100100000" OR uut_h_0_1 /= "111111111111100110100110101110" OR uut_h_0_2 /= "111111110000010101011000111111" OR uut_h_1_0 /= "000000000001010101010111100001" OR uut_h_1_1 /= "000000000000001101111000111010" OR uut_h_1_2 /= "111111111101100110111111000111" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "000010";
              state <= "111110";
            ELSE
              state <= "000110";
            END IF;
            uut_rst <= '0';
          WHEN "000110" =>
            uut_h_0_0_i <= "000000001100011011110010001";
            uut_h_0_1_i <= "000000001010110111100111100";
            uut_h_0_2_i <= "111111110111011000100111001";
            uut_h_1_0_i <= "111111111000011011111111001";
            uut_h_1_1_i <= "111111111111110110110111011";
            uut_h_1_2_i <= "000000000101000011011111010";
            uut_coord_trans <= "111111010110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111110001001100010100000" OR uut_h_0_1 /= "000000000001101000110111011000" OR uut_h_0_2 /= "111111100111110010100001111001" OR uut_h_1_0 /= "000000000001111001110011011110" OR uut_h_1_1 /= "111111111111100010000111001000" OR uut_h_1_2 /= "111111111011101101110101000110" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "000011";
              state <= "111110";
            ELSE
              state <= "000111";
            END IF;
            uut_rst <= '0';
          WHEN "000111" =>
            uut_h_0_0_i <= "000000000011111010011110110";
            uut_h_0_1_i <= "111111111101001100010101011";
            uut_h_0_2_i <= "111111110100010101011110100";
            uut_h_1_0_i <= "000000000110111010001011001";
            uut_h_1_1_i <= "111111111011100101110011000";
            uut_h_1_2_i <= "000000001100110111011100000";
            uut_coord_trans <= "111111111111";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000100000000000010100" OR uut_h_0_1 /= "111111111110110110110100111001" OR uut_h_0_2 /= "111111001010000100110100010010" OR uut_h_1_0 /= "000000000000010001010011100000" OR uut_h_1_1 /= "111111111110000000111111001110" OR uut_h_1_2 /= "111110110100101100100010001111" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "000100";
              state <= "111110";
            ELSE
              state <= "001000";
            END IF;
            uut_rst <= '0';
          WHEN "001000" =>
            uut_h_0_0_i <= "000000001001000100110010110";
            uut_h_0_1_i <= "000000000110010010101011010";
            uut_h_0_2_i <= "000000001100010111010111110";
            uut_h_1_0_i <= "000000000101101010100111111";
            uut_h_1_1_i <= "111111110100001000001101111";
            uut_h_1_2_i <= "000000000000011110101110101";
            uut_coord_trans <= "000001011111";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000001010011010110111110" OR uut_h_0_1 /= "111111111111100100000010110010" OR uut_h_0_2 /= "000000000011111001110101011101" OR uut_h_1_0 /= "000000000001100010001110010110" OR uut_h_1_1 /= "000000000001001101001000110100" OR uut_h_1_2 /= "111111111110100100110110101101" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "000101";
              state <= "111110";
            ELSE
              state <= "001001";
            END IF;
            uut_rst <= '0';
          WHEN "001001" =>
            uut_h_0_0_i <= "111111110100000000111100010";
            uut_h_0_1_i <= "000000001001000000010111101";
            uut_h_0_2_i <= "111111110000011101100110110";
            uut_h_1_0_i <= "000000001000000100100110000";
            uut_h_1_1_i <= "111111110110000110111011010";
            uut_h_1_2_i <= "111111111010011010001011110";
            uut_coord_trans <= "111111110110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000001100011011110010001" OR uut_h_0_1 /= "000000000001010110111100111100" OR uut_h_0_2 /= "000000010010000110000000001010" OR uut_h_1_0 /= "111111111111000011011111111001" OR uut_h_1_1 /= "111111111111111110110110111011" OR uut_h_1_2 /= "111111000010011001111010111110" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "000110";
              state <= "111110";
            ELSE
              state <= "001010";
            END IF;
            uut_rst <= '0';
          WHEN "001010" =>
            uut_h_0_0_i <= "000000000010010100000001001";
            uut_h_0_1_i <= "000000000001000010101000101";
            uut_h_0_2_i <= "000000000001011011110100011";
            uut_h_1_0_i <= "000000001001010110000100000";
            uut_h_1_1_i <= "000000001101100111110101111";
            uut_h_1_2_i <= "000000001100110101100000000";
            uut_coord_trans <= "000000111101";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000011111010011110110" OR uut_h_0_1 /= "111111111111101001100010101011" OR uut_h_0_2 /= "111111111101100111000111000101" OR uut_h_1_0 /= "000000000000110111010001011001" OR uut_h_1_1 /= "111111111111011100101110011000" OR uut_h_1_2 /= "000000000000110000111011011001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "000111";
              state <= "111110";
            ELSE
              state <= "001011";
            END IF;
            uut_rst <= '0';
          WHEN "001011" =>
            uut_h_0_0_i <= "111111111010101101111000100";
            uut_h_0_1_i <= "111111111011001001001011110";
            uut_h_0_2_i <= "000000001110100100100110001";
            uut_h_1_0_i <= "111111110111010100010101111";
            uut_h_1_1_i <= "111111110101010010111000100";
            uut_h_1_2_i <= "000000000101110001001111000";
            uut_coord_trans <= "000001010111";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000001001000100110010110" OR uut_h_0_1 /= "000000000000110010010101011010" OR uut_h_0_2 /= "000000000101010011100100110110" OR uut_h_1_0 /= "000000000000101101010100111111" OR uut_h_1_1 /= "111111111110100001000001101111" OR uut_h_1_2 /= "000010000011111001111110101101" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "001000";
              state <= "111110";
            ELSE
              state <= "001100";
            END IF;
            uut_rst <= '0';
          WHEN "001100" =>
            uut_h_0_0_i <= "000000000101110001000010011";
            uut_h_0_1_i <= "000000001100010101101111101";
            uut_h_0_2_i <= "111111110010010110010011011";
            uut_h_1_0_i <= "000000001101010110111000100";
            uut_h_1_1_i <= "000000001101011100001111110";
            uut_h_1_2_i <= "000000001000100011101000011";
            uut_coord_trans <= "000000101101";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111110100000000111100010" OR uut_h_0_1 /= "000000000001001000000010111101" OR uut_h_0_2 /= "111111110010001100100001010001" OR uut_h_1_0 /= "000000000001000000100100110000" OR uut_h_1_1 /= "111111111110110000110111011010" OR uut_h_1_2 /= "111111110100001010011110010000" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "001001";
              state <= "111110";
            ELSE
              state <= "001101";
            END IF;
            uut_rst <= '0';
          WHEN "001101" =>
            uut_h_0_0_i <= "111111111110010101010001110";
            uut_h_0_1_i <= "000000000001000000011010000";
            uut_h_0_2_i <= "111111111111000011010100100";
            uut_h_1_0_i <= "000000000100110101110000011";
            uut_h_1_1_i <= "000000000100010010000001100";
            uut_h_1_2_i <= "000000001100010111001100100";
            uut_coord_trans <= "111111110100";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000010010100000001001" OR uut_h_0_1 /= "000000000000001000010101000101" OR uut_h_0_2 /= "000000110000011001000111011001" OR uut_h_1_0 /= "000000000001001010110000100000" OR uut_h_1_1 /= "000000000001101100111110101111" OR uut_h_1_2 /= "111111100111000010101011010111" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "001010";
              state <= "111110";
            ELSE
              state <= "001110";
            END IF;
            uut_rst <= '0';
          WHEN "001110" =>
            uut_h_0_0_i <= "000000000101000110110000010";
            uut_h_0_1_i <= "000000000110001101111001011";
            uut_h_0_2_i <= "000000001100001000110000110";
            uut_h_1_0_i <= "111111111001011011101100011";
            uut_h_1_1_i <= "111111110110100111100010100";
            uut_h_1_2_i <= "000000000001110110011111100";
            uut_coord_trans <= "000001001110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111111010101101111000100" OR uut_h_0_1 /= "111111111111011001001001011110" OR uut_h_0_2 /= "000010001111111101001001101010" OR uut_h_1_0 /= "111111111110111010100010101111" OR uut_h_1_1 /= "111111111110101010010111000100" OR uut_h_1_2 /= "000011000001001000110111101110" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "001011";
              state <= "111110";
            ELSE
              state <= "001111";
            END IF;
            uut_rst <= '0';
          WHEN "001111" =>
            uut_h_0_0_i <= "000000001010111100000110001";
            uut_h_0_1_i <= "111111110100111010101001111";
            uut_h_0_2_i <= "000000000011000101100010000";
            uut_h_1_0_i <= "111111110100001011111111101";
            uut_h_1_1_i <= "111111110000111011001100010";
            uut_h_1_2_i <= "000000000011011111010101010";
            uut_coord_trans <= "000000101110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000101110001000010011" OR uut_h_0_1 /= "000000000001100010101101111101" OR uut_h_0_2 /= "111111111000010111101101110100" OR uut_h_1_0 /= "000000000001101010110111000100" OR uut_h_1_1 /= "000000000001101011100001111110" OR uut_h_1_2 /= "111111100010101100101001110110" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "001100";
              state <= "111110";
            ELSE
              state <= "010000";
            END IF;
            uut_rst <= '0';
          WHEN "010000" =>
            uut_h_0_0_i <= "111111111001101000101111111";
            uut_h_0_1_i <= "000000000111011100111000101";
            uut_h_0_2_i <= "000000001001111010011100101";
            uut_h_1_0_i <= "111111111111110110111011111";
            uut_h_1_1_i <= "111111110011101111001000000";
            uut_h_1_2_i <= "000000000111110110001111010";
            uut_coord_trans <= "000000010000";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111111110010101010001110" OR uut_h_0_1 /= "000000000000001000000011010000" OR uut_h_0_2 /= "111111110011011000101011011000" OR uut_h_1_0 /= "000000000000100110101110000011" OR uut_h_1_1 /= "000000000000100010010000001100" OR uut_h_1_2 /= "111111111100011000101110111110" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "001101";
              state <= "111110";
            ELSE
              state <= "010001";
            END IF;
            uut_rst <= '0';
          WHEN "010001" =>
            uut_h_0_0_i <= "111111111111000000011010011";
            uut_h_0_1_i <= "000000000101111100110100001";
            uut_h_0_2_i <= "111111110101111000010111101";
            uut_h_1_0_i <= "111111110010110010101110000";
            uut_h_1_1_i <= "111111111000100011011110110";
            uut_h_1_2_i <= "111111111001100110010001110";
            uut_coord_trans <= "111111001011";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000101000110110000010" OR uut_h_0_1 /= "000000000000110001101111001011" OR uut_h_0_2 /= "000000011000010100011011001011" OR uut_h_1_0 /= "111111111111001011011101100011" OR uut_h_1_1 /= "111111111110110100111100010100" OR uut_h_1_2 /= "000010011011111111000011011011" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "001110";
              state <= "111110";
            ELSE
              state <= "010010";
            END IF;
            uut_rst <= '0';
          WHEN "010010" =>
            uut_h_0_0_i <= "111111110110001111011110010";
            uut_h_0_1_i <= "000000000000101101101111001";
            uut_h_0_2_i <= "000000001101100110111000000";
            uut_h_1_0_i <= "000000000110100100100111011";
            uut_h_1_1_i <= "111111111001011110100011110";
            uut_h_1_2_i <= "111111110110111010001001000";
            uut_coord_trans <= "000001010001";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000001010111100000110001" OR uut_h_0_1 /= "111111111110100111010101001111" OR uut_h_0_2 /= "000000101110110011010010010000" OR uut_h_1_0 /= "111111111110100001011111111101" OR uut_h_1_1 /= "111111111110000111011001100010" OR uut_h_1_2 /= "000001111011101111010000100001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "001111";
              state <= "111110";
            ELSE
              state <= "010011";
            END IF;
            uut_rst <= '0';
          WHEN "010011" =>
            uut_h_0_0_i <= "000000000101110000101110011";
            uut_h_0_1_i <= "111111110011010010110001101";
            uut_h_0_2_i <= "000000000100000000011111110";
            uut_h_1_0_i <= "000000000000011110100111110";
            uut_h_1_1_i <= "000000001111111001100111000";
            uut_h_1_2_i <= "111111111100100101100111010";
            uut_coord_trans <= "000000001001";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111111001101000101111111" OR uut_h_0_1 /= "000000000000111011100111000101" OR uut_h_0_2 /= "000000010000001001101011000101" OR uut_h_1_0 /= "111111111111111110110111011111" OR uut_h_1_1 /= "111111111110011101111001000000" OR uut_h_1_2 /= "000000011101011000101110000010" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "010000";
              state <= "111110";
            ELSE
              state <= "010100";
            END IF;
            uut_rst <= '0';
          WHEN "010100" =>
            uut_h_0_0_i <= "000000000000010010101010000";
            uut_h_0_1_i <= "000000001010111011110111001";
            uut_h_0_2_i <= "000000001001000100011100010";
            uut_h_1_0_i <= "111111110111111001011001110";
            uut_h_1_1_i <= "111111110001100010110100001";
            uut_h_1_2_i <= "000000001111000111011110011";
            uut_coord_trans <= "000000110111";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111111111000000011010011" OR uut_h_0_1 /= "000000000000101111100110100001" OR uut_h_0_2 /= "111111011010001001110111000000" OR uut_h_1_0 /= "111111111110010110010101110000" OR uut_h_1_1 /= "111111111111000100011011110110" OR uut_h_1_2 /= "111110000101110010010100011101" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "010001";
              state <= "111110";
            ELSE
              state <= "010101";
            END IF;
            uut_rst <= '0';
          WHEN "010101" =>
            uut_h_0_0_i <= "000000000111010010010100110";
            uut_h_0_1_i <= "000000001110000010100111101";
            uut_h_0_2_i <= "000000000101011101000110001";
            uut_h_1_0_i <= "000000000100110101001110001";
            uut_h_1_1_i <= "000000000001000111110110001";
            uut_h_1_2_i <= "111111111110000110001101101";
            uut_coord_trans <= "111111110011";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111110110001111011110010" OR uut_h_0_1 /= "000000000000000101101101111001" OR uut_h_0_2 /= "000010000000011110111111010011" OR uut_h_1_0 /= "000000000000110100100100111011" OR uut_h_1_1 /= "111111111111001011110100011110" OR uut_h_1_2 /= "000001001111100111001100110100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "010010";
              state <= "111110";
            ELSE
              state <= "010110";
            END IF;
            uut_rst <= '0';
          WHEN "010110" =>
            uut_h_0_0_i <= "000000000001100001100100101";
            uut_h_0_1_i <= "000000001000000010110000110";
            uut_h_0_2_i <= "111111110010110101100111010";
            uut_h_1_0_i <= "111111111100101001001111010";
            uut_h_1_1_i <= "000000000000101101110001100";
            uut_h_1_2_i <= "111111111000000001101111101";
            uut_coord_trans <= "000000011011";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000101110000101110011" OR uut_h_0_1 /= "111111111110011010010110001101" OR uut_h_0_2 /= "000000001101011010000101111111" OR uut_h_1_0 /= "000000000000000011110100111110" OR uut_h_1_1 /= "000000000001111111001100111000" OR uut_h_1_2 /= "111111111111010111000100100111" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "010011";
              state <= "111110";
            ELSE
              state <= "010111";
            END IF;
            uut_rst <= '0';
          WHEN "010111" =>
            uut_h_0_0_i <= "000000000110101100111100011";
            uut_h_0_1_i <= "111111110010111100111000101";
            uut_h_0_2_i <= "000000001111000011011111011";
            uut_h_1_0_i <= "000000001111110000111000101";
            uut_h_1_1_i <= "000000001110100000110110011";
            uut_h_1_2_i <= "000000000011000110101010110";
            uut_coord_trans <= "111110101010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000000010010101010000" OR uut_h_0_1 /= "000000000001010111011110111001" OR uut_h_0_2 /= "000000010001100010101001101011" OR uut_h_1_0 /= "111111111110111111001011001110" OR uut_h_1_1 /= "111111111110001100010110100001" OR uut_h_1_2 /= "000010000110011011111100000111" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "010100";
              state <= "111110";
            ELSE
              state <= "011000";
            END IF;
            uut_rst <= '0';
          WHEN "011000" =>
            uut_h_0_0_i <= "111111111001100110011111000";
            uut_h_0_1_i <= "111111111011010101111101011";
            uut_h_0_2_i <= "111111110001111111010001101";
            uut_h_1_0_i <= "000000001010000010001000111";
            uut_h_1_1_i <= "111111110100001110010110111";
            uut_h_1_2_i <= "000000000110011101011000000";
            uut_coord_trans <= "000000010111";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000111010010010100110" OR uut_h_0_1 /= "000000000001110000010100111101" OR uut_h_0_2 /= "000000000101000000101001110101" OR uut_h_1_0 /= "000000000000100110101001110001" OR uut_h_1_1 /= "000000000000001000111110110001" OR uut_h_1_2 /= "111111110111100110011001001011" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "010101";
              state <= "111110";
            ELSE
              state <= "011001";
            END IF;
            uut_rst <= '0';
          WHEN "011001" =>
            uut_h_0_0_i <= "111111110101100011111000100";
            uut_h_0_1_i <= "111111111001000110101011011";
            uut_h_0_2_i <= "000000001110000001010111101";
            uut_h_1_0_i <= "000000000100110110000100011";
            uut_h_1_1_i <= "000000001010100100111111001";
            uut_h_1_2_i <= "111111110000000000101010101";
            uut_coord_trans <= "111110011101";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000001100001100100101" OR uut_h_0_1 /= "000000000001000000010110000110" OR uut_h_0_2 /= "000000001001001101011000110110" OR uut_h_1_0 /= "111111111111100101001001111010" OR uut_h_1_1 /= "000000000000000101101110001100" OR uut_h_1_2 /= "000000011110011101011000101100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "010110";
              state <= "111110";
            ELSE
              state <= "011010";
            END IF;
            uut_rst <= '0';
          WHEN "011010" =>
            uut_h_0_0_i <= "111111110011011001111100110";
            uut_h_0_1_i <= "111111110111101010101101110";
            uut_h_0_2_i <= "111111111100011000101101010";
            uut_h_1_0_i <= "111111110011011010101101110";
            uut_h_1_1_i <= "111111111011000100111001010";
            uut_h_1_2_i <= "111111111101011110010010010";
            uut_coord_trans <= "000000111001";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000110101100111100011" OR uut_h_0_1 /= "111111111110010111100111000101" OR uut_h_0_2 /= "111110001001110001010000110011" OR uut_h_1_0 /= "000000000001111110000111000101" OR uut_h_1_1 /= "000000000001110100000110110011" OR uut_h_1_2 /= "000001001101001000001001111110" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "010111";
              state <= "111110";
            ELSE
              state <= "011011";
            END IF;
            uut_rst <= '0';
          WHEN "011011" =>
            uut_h_0_0_i <= "111111111000101000111100101";
            uut_h_0_1_i <= "000000001010011011110110110";
            uut_h_0_2_i <= "000000000011100001111111110";
            uut_h_1_0_i <= "000000001011000000011110011";
            uut_h_1_1_i <= "111111110101110101001000010";
            uut_h_1_2_i <= "000000000110011100110001111";
            uut_coord_trans <= "111110101111";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111111001100110011111000" OR uut_h_0_1 /= "111111111111011010101111101011" OR uut_h_0_2 /= "000000100101001001000001011011" OR uut_h_1_0 /= "000000000001010000010001000111" OR uut_h_1_1 /= "111111111110100001110010110111" OR uut_h_1_2 /= "000000011010010011111101011000" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "011000";
              state <= "111110";
            ELSE
              state <= "011100";
            END IF;
            uut_rst <= '0';
          WHEN "011100" =>
            uut_h_0_0_i <= "000000000011001000010111010";
            uut_h_0_1_i <= "111111110010110111001010101";
            uut_h_0_2_i <= "111111111110011110001010111";
            uut_h_1_0_i <= "000000001001111111011100111";
            uut_h_1_1_i <= "000000000111011001101010001";
            uut_h_1_2_i <= "111111110010010000110001001";
            uut_coord_trans <= "000000101110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111110101100011111000100" OR uut_h_0_1 /= "111111111111001000110101011011" OR uut_h_0_2 /= "111100110011011111100000111100" OR uut_h_1_0 /= "000000000000100110110000100011" OR uut_h_1_1 /= "000000000001010100100111111001" OR uut_h_1_2 /= "111111111010011011011111000000" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "011001";
              state <= "111110";
            ELSE
              state <= "011101";
            END IF;
            uut_rst <= '0';
          WHEN "011101" =>
            uut_h_0_0_i <= "111111110001010010111011010";
            uut_h_0_1_i <= "000000001110100001011100000";
            uut_h_0_2_i <= "000000000100101011011101010";
            uut_h_1_0_i <= "111111111101100101011011000";
            uut_h_1_1_i <= "111111110110101011110101101";
            uut_h_1_2_i <= "111111110011011110000001101";
            uut_coord_trans <= "111111001101";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111110011011001111100110" OR uut_h_0_1 /= "111111111110111101010101101110" OR uut_h_0_2 /= "000010000011000110011110010000" OR uut_h_1_0 /= "111111111110011011010101101110" OR uut_h_1_1 /= "111111111111011000100111001010" OR uut_h_1_2 /= "000001110111000011001011010110" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "011010";
              state <= "111110";
            ELSE
              state <= "011110";
            END IF;
            uut_rst <= '0';
          WHEN "011110" =>
            uut_h_0_0_i <= "000000000011011001110100010";
            uut_h_0_1_i <= "111111111111101001100011010";
            uut_h_0_2_i <= "000000001100110101001100100";
            uut_h_1_0_i <= "000000001010001000100101111";
            uut_h_1_1_i <= "000000001000010101111110001";
            uut_h_1_2_i <= "111111110110110110110000100";
            uut_coord_trans <= "000000111000";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111111000101000111100101" OR uut_h_0_1 /= "000000000001010011011110110110" OR uut_h_0_2 /= "111110111111000000100100000100" OR uut_h_1_0 /= "000000000001011000000011110011" OR uut_h_1_1 /= "111111111110101110101001000010" OR uut_h_1_2 /= "111110110100000010111101110010" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "011011";
              state <= "111110";
            ELSE
              state <= "011111";
            END IF;
            uut_rst <= '0';
          WHEN "011111" =>
            uut_h_0_0_i <= "111111110110001110001101110";
            uut_h_0_1_i <= "000000000010101010100000110";
            uut_h_0_2_i <= "111111111001100010100100110";
            uut_h_1_0_i <= "000000000111111001101000010";
            uut_h_1_1_i <= "111111111000010101100110100";
            uut_h_1_2_i <= "000000001101010110010001111";
            uut_coord_trans <= "111111010001";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000011001000010111010" OR uut_h_0_1 /= "111111111110010110111001010101" OR uut_h_0_2 /= "000001001010100101000111111110" OR uut_h_1_0 /= "000000000001001111111011100111" OR uut_h_1_1 /= "000000000000111011001101010001" OR uut_h_1_2 /= "111111111010010001111010000001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "011100";
              state <= "111110";
            ELSE
              state <= "100000";
            END IF;
            uut_rst <= '0';
          WHEN "100000" =>
            uut_h_0_0_i <= "000000001000011010100100000";
            uut_h_0_1_i <= "000000001100001010001101100";
            uut_h_0_2_i <= "000000000101011010001100111";
            uut_h_1_0_i <= "000000001000101101011010001";
            uut_h_1_1_i <= "000000001001100010101001110";
            uut_h_1_2_i <= "111111111001011110110011110";
            uut_coord_trans <= "111111010100";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111110001010010111011010" OR uut_h_0_1 /= "000000000001110100001011100000" OR uut_h_0_2 /= "111111001101000000010101110001" OR uut_h_1_0 /= "111111111111101100101011011000" OR uut_h_1_1 /= "111111111110110101011110101101" OR uut_h_1_2 /= "111110100110000010110001001101" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "011101";
              state <= "111110";
            ELSE
              state <= "100001";
            END IF;
            uut_rst <= '0';
          WHEN "100001" =>
            uut_h_0_0_i <= "111111110101011001110111011";
            uut_h_0_1_i <= "000000000100111010010000010";
            uut_h_0_2_i <= "111111110010011100100011000";
            uut_h_1_0_i <= "000000000111110110000110011";
            uut_h_1_1_i <= "000000001110111011100011000";
            uut_h_1_2_i <= "000000001001010100110100010";
            uut_coord_trans <= "000000010001";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000011011001110100010" OR uut_h_0_1 /= "111111111111111101001100011010" OR uut_h_0_2 /= "000000101110111010110111010100" OR uut_h_1_0 /= "000000000001010001000100101111" OR uut_h_1_1 /= "000000000001000010101111110001" OR uut_h_1_2 /= "111111110110001011111000000100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "011110";
              state <= "111110";
            ELSE
              state <= "100010";
            END IF;
            uut_rst <= '0';
          WHEN "100010" =>
            uut_h_0_0_i <= "111111110101110111011110010";
            uut_h_0_1_i <= "000000001010011101011100010";
            uut_h_0_2_i <= "000000000100110100101110111";
            uut_h_1_0_i <= "111111110010011101100001111";
            uut_h_1_1_i <= "111111111001101000010111000";
            uut_h_1_2_i <= "000000001010001001111110011";
            uut_coord_trans <= "111111100110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111110110001110001101110" OR uut_h_0_1 /= "000000000000010101010100000110" OR uut_h_0_2 /= "111110111011010010111101001100" OR uut_h_1_0 /= "000000000000111111001101000010" OR uut_h_1_1 /= "111111111111000010101100110100" OR uut_h_1_2 /= "111111010011010111100001100100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "011111";
              state <= "111110";
            ELSE
              state <= "100011";
            END IF;
            uut_rst <= '0';
          WHEN "100011" =>
            uut_h_0_0_i <= "111111110110000100110101101";
            uut_h_0_1_i <= "111111111001000011010110101";
            uut_h_0_2_i <= "111111111010011010001100010";
            uut_h_1_0_i <= "000000000100101100000010010";
            uut_h_1_1_i <= "000000000100011011110110101";
            uut_h_1_2_i <= "000000001111101001010111110";
            uut_coord_trans <= "000000101111";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000001000011010100100000" OR uut_h_0_1 /= "000000000001100001010001101100" OR uut_h_0_2 /= "000000001101010000011001101111" OR uut_h_1_0 /= "000000000001000101101011010001" OR uut_h_1_1 /= "000000000001001100010101001110" OR uut_h_1_2 /= "000000000101011000000001001000" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "100000";
              state <= "111110";
            ELSE
              state <= "100100";
            END IF;
            uut_rst <= '0';
          WHEN "100100" =>
            uut_h_0_0_i <= "111111110101000000110000000";
            uut_h_0_1_i <= "111111111011100001000110000";
            uut_h_0_2_i <= "111111111000110001000000100";
            uut_h_1_0_i <= "111111111101111010001010000";
            uut_h_1_1_i <= "111111110010011100001000101";
            uut_h_1_2_i <= "111111110100001110011100101";
            uut_coord_trans <= "111111111101";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111110101011001110111011" OR uut_h_0_1 /= "000000000000100111010010000010" OR uut_h_0_2 /= "000000010101010110001100010010" OR uut_h_1_0 /= "000000000000111110110000110011" OR uut_h_1_1 /= "000000000001110111011100011000" OR uut_h_1_2 /= "111111111001111101110110100101" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "100001";
              state <= "111110";
            ELSE
              state <= "100101";
            END IF;
            uut_rst <= '0';
          WHEN "100101" =>
            uut_h_0_0_i <= "111111110011110011101010010";
            uut_h_0_1_i <= "000000001100010001101001001";
            uut_h_0_2_i <= "111111110010010000111011000";
            uut_h_1_0_i <= "000000001101101001100010011";
            uut_h_1_1_i <= "111111111101100101010100111";
            uut_h_1_2_i <= "000000001101100101111011110";
            uut_coord_trans <= "111110110000";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111110101110111011110010" OR uut_h_0_1 /= "000000000001010011101011100010" OR uut_h_0_2 /= "111111100111001000100100111011" OR uut_h_1_0 /= "111111111110010011101100001111" OR uut_h_1_1 /= "111111111111001101000010111000" OR uut_h_1_2 /= "111111000110111010110100001110" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "100010";
              state <= "111110";
            ELSE
              state <= "100110";
            END IF;
            uut_rst <= '0';
          WHEN "100110" =>
            uut_h_0_0_i <= "000000000110011010000011111";
            uut_h_0_1_i <= "111111110110110111010000001";
            uut_h_0_2_i <= "000000000110011111110000001";
            uut_h_1_0_i <= "111111111100101010100110110";
            uut_h_1_1_i <= "111111110111111101100010100";
            uut_h_1_2_i <= "000000001000001000100000010";
            uut_coord_trans <= "000000001010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111110110000100110101101" OR uut_h_0_1 /= "111111111111001000011010110101" OR uut_h_0_2 /= "000001011111110111001101100100" OR uut_h_1_0 /= "000000000000100101100000010010" OR uut_h_1_1 /= "000000000000100011011110110101" OR uut_h_1_2 /= "000000010110001001111111111010" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "100011";
              state <= "111110";
            ELSE
              state <= "100111";
            END IF;
            uut_rst <= '0';
          WHEN "100111" =>
            uut_h_0_0_i <= "000000000100001011011010011";
            uut_h_0_1_i <= "000000000011001101101110111";
            uut_h_0_2_i <= "111111111010101110111100001";
            uut_h_1_0_i <= "000000001111100010001101110";
            uut_h_1_1_i <= "000000001101000110000000111";
            uut_h_1_2_i <= "000000001110101000001110001";
            uut_coord_trans <= "000000010100";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111110101000000110000000" OR uut_h_0_1 /= "111111111111011100001000110000" OR uut_h_0_2 /= "111111111001001100011110001100" OR uut_h_1_0 /= "111111111111101111010001010000" OR uut_h_1_1 /= "111111111110010011100001000101" OR uut_h_1_2 /= "111111111000100101111111000101" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "100100";
              state <= "111110";
            ELSE
              state <= "101000";
            END IF;
            uut_rst <= '0';
          WHEN "101000" =>
            uut_h_0_0_i <= "000000000111000011000110001";
            uut_h_0_1_i <= "111111110010100111001010100";
            uut_h_0_2_i <= "000000000001111001100100000";
            uut_h_1_0_i <= "000000000101101110001000110";
            uut_h_1_1_i <= "111111111000110010001000100";
            uut_h_1_2_i <= "111111111110110111100011101";
            uut_coord_trans <= "000000110110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111110011110011101010010" OR uut_h_0_1 /= "000000000001100010001101001001" OR uut_h_0_2 /= "111110101110101100101000010000" OR uut_h_1_0 /= "000000000001101101001100010011" OR uut_h_1_1 /= "111111111111101100101010100111" OR uut_h_1_2 /= "111111101001110111000011101110" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "100101";
              state <= "111110";
            ELSE
              state <= "101001";
            END IF;
            uut_rst <= '0';
          WHEN "101001" =>
            uut_h_0_0_i <= "000000000100111011001110101";
            uut_h_0_1_i <= "111111111101110101100000011";
            uut_h_0_2_i <= "111111111111010111110011010";
            uut_h_1_0_i <= "000000000101000011000001111";
            uut_h_1_1_i <= "000000000000001010011010101";
            uut_h_1_2_i <= "111111111010111101010001110";
            uut_coord_trans <= "111111101000";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000110011010000011111" OR uut_h_0_1 /= "111111111110110110111010000001" OR uut_h_0_2 /= "000000001100100001001001100001" OR uut_h_1_0 /= "111111111111100101010100110110" OR uut_h_1_1 /= "111111111110111111101100010100" OR uut_h_1_2 /= "000000010010000111111110010000" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "100110";
              state <= "111110";
            ELSE
              state <= "101010";
            END IF;
            uut_rst <= '0';
          WHEN "101010" =>
            uut_h_0_0_i <= "000000000110110001010001000";
            uut_h_0_1_i <= "000000001110000000000111110";
            uut_h_0_2_i <= "111111110110111110110110111";
            uut_h_1_0_i <= "111111111111011000111100111";
            uut_h_1_1_i <= "000000000000100011010101100";
            uut_h_1_2_i <= "000000001011111100010110100";
            uut_coord_trans <= "111111111001";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000100001011011010011" OR uut_h_0_1 /= "000000000000011001101101110111" OR uut_h_0_2 /= "000000001010000110011011111101" OR uut_h_1_0 /= "000000000001111100010001101110" OR uut_h_1_1 /= "000000000001101000110000000111" OR uut_h_1_2 /= "111111110010000010101111011111" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "100111";
              state <= "111110";
            ELSE
              state <= "101011";
            END IF;
            uut_rst <= '0';
          WHEN "101011" =>
            uut_h_0_0_i <= "111111110000101100111010011";
            uut_h_0_1_i <= "111111110101010010101110010";
            uut_h_0_2_i <= "111111110110110101110010011";
            uut_h_1_0_i <= "000000001001110111010110111";
            uut_h_1_1_i <= "111111110101110011111011001";
            uut_h_1_2_i <= "111111111001100010100001001";
            uut_coord_trans <= "000000000000";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000111000011000110001" OR uut_h_0_1 /= "111111111110010100111001010100" OR uut_h_0_2 /= "000001001011101000100100011001" OR uut_h_1_0 /= "000000000000101101110001000110" OR uut_h_1_1 /= "111111111111000110010001000100" OR uut_h_1_2 /= "000000111010111010000010001111" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "101000";
              state <= "111110";
            ELSE
              state <= "101100";
            END IF;
            uut_rst <= '0';
          WHEN "101100" =>
            uut_h_0_0_i <= "000000001101000110100101010";
            uut_h_0_1_i <= "000000000010010011111110100";
            uut_h_0_2_i <= "111111110100000010010000000";
            uut_h_1_0_i <= "111111110001110110011110111";
            uut_h_1_1_i <= "000000000010000101010000011";
            uut_h_1_2_i <= "111111111001100110101000111";
            uut_coord_trans <= "000001011010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000100111011001110101" OR uut_h_0_1 /= "111111111111101110101100000011" OR uut_h_0_2 /= "111111101100000100000100111010" OR uut_h_1_0 /= "000000000000101000011000001111" OR uut_h_1_1 /= "000000000000000001010011010101" OR uut_h_1_2 /= "111111101111001011110100111110" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "101001";
              state <= "111110";
            ELSE
              state <= "101101";
            END IF;
            uut_rst <= '0';
          WHEN "101101" =>
            uut_h_0_0_i <= "000000001000100001011000011";
            uut_h_0_1_i <= "111111111011001011011010000";
            uut_h_0_2_i <= "000000001001111000000111101";
            uut_h_1_0_i <= "000000001000000010101010111";
            uut_h_1_1_i <= "111111110100110101111100100";
            uut_h_1_2_i <= "000000000100010000000111011";
            uut_coord_trans <= "000000011011";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000110110001010001000" OR uut_h_0_1 /= "000000000001110000000000111110" OR uut_h_0_2 /= "000000000000111101011101101100" OR uut_h_1_0 /= "111111111111111011000111100111" OR uut_h_1_1 /= "000000000000000100011010101100" OR uut_h_1_2 /= "111111111010011101111010110111" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "101010";
              state <= "111110";
            ELSE
              state <= "101110";
            END IF;
            uut_rst <= '0';
          WHEN "101110" =>
            uut_h_0_0_i <= "000000000111010101101001101";
            uut_h_0_1_i <= "111111110101110001110110011";
            uut_h_0_2_i <= "000000001100111111100110000";
            uut_h_1_0_i <= "000000001011100000111101101";
            uut_h_1_1_i <= "000000000010010110001000011";
            uut_h_1_2_i <= "111111110010011110011001011";
            uut_coord_trans <= "000000010000";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111110000101100111010011" OR uut_h_0_1 /= "111111111110101010010101110010" OR uut_h_0_2 /= "111111111110110110101110010011" OR uut_h_1_0 /= "000000000001001110111010110111" OR uut_h_1_1 /= "111111111110101110011111011001" OR uut_h_1_2 /= "111111111111001100010100001001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "101011";
              state <= "111110";
            ELSE
              state <= "101111";
            END IF;
            uut_rst <= '0';
          WHEN "101111" =>
            uut_h_0_0_i <= "111111111111001101010010000";
            uut_h_0_1_i <= "111111110111010001100010000";
            uut_h_0_2_i <= "000000000101000011110100100";
            uut_h_1_0_i <= "000000001001110001010010111";
            uut_h_1_1_i <= "000000000110101101000001100";
            uut_h_1_2_i <= "000000000100010010011001010";
            uut_coord_trans <= "111111000000";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000001101000110100101010" OR uut_h_0_1 /= "000000000000010010011111110100" OR uut_h_0_2 /= "000000000001110010111000111010" OR uut_h_1_0 /= "111111111110001110110011110111" OR uut_h_1_1 /= "000000000000010000101010000011" OR uut_h_1_2 /= "000010011101000100110011010101" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "101100";
              state <= "111110";
            ELSE
              state <= "110000";
            END IF;
            uut_rst <= '0';
          WHEN "110000" =>
            uut_h_0_0_i <= "111111110101010100101100001";
            uut_h_0_1_i <= "000000001110100011110000010";
            uut_h_0_2_i <= "111111110000110100100111100";
            uut_h_1_0_i <= "111111110100110010011001010";
            uut_h_1_1_i <= "111111110000100000100101001";
            uut_h_1_2_i <= "000000001111000100110101011";
            uut_coord_trans <= "000000000101";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000001000100001011000011" OR uut_h_0_1 /= "111111111111011001011011010000" OR uut_h_0_2 /= "000000010101111111011011111101" OR uut_h_1_0 /= "000000000001000000010101010111" OR uut_h_1_1 /= "111111111110100110101111100100" OR uut_h_1_2 /= "000000100000110010011110011111" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "101101";
              state <= "111110";
            ELSE
              state <= "110001";
            END IF;
            uut_rst <= '0';
          WHEN "110001" =>
            uut_h_0_0_i <= "000000001011100110000100100";
            uut_h_0_1_i <= "000000000101001001001001110";
            uut_h_0_2_i <= "111111110011011101000011010";
            uut_h_1_0_i <= "000000001100101011110101100";
            uut_h_1_1_i <= "000000001110000111101001000";
            uut_h_1_2_i <= "111111110101101110011000101";
            uut_coord_trans <= "111110100101";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000111010101101001101" OR uut_h_0_1 /= "111111111110101110001110110011" OR uut_h_0_2 /= "000000010100100000011100110000" OR uut_h_1_0 /= "000000000001011100000111101101" OR uut_h_1_1 /= "000000000000010010110001000011" OR uut_h_1_2 /= "000000000000011100101101001011" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "101110";
              state <= "111110";
            ELSE
              state <= "110010";
            END IF;
            uut_rst <= '0';
          WHEN "110010" =>
            uut_h_0_0_i <= "111111110010010001111111011";
            uut_h_0_1_i <= "000000001111111001111100001";
            uut_h_0_2_i <= "000000001011100100000010101";
            uut_h_1_0_i <= "111111111111101001101110101";
            uut_h_1_1_i <= "111111110000001000111111101";
            uut_h_1_2_i <= "000000001101000101111010101";
            uut_coord_trans <= "000001001011";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111111111001101010010000" OR uut_h_0_1 /= "111111111110111010001100010000" OR uut_h_0_2 /= "111110011010100011101110100100" OR uut_h_1_0 /= "000000000001001110001010010111" OR uut_h_1_1 /= "000000000000110101101000001100" OR uut_h_1_2 /= "000000000010011011100100101010" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "101111";
              state <= "111110";
            ELSE
              state <= "110011";
            END IF;
            uut_rst <= '0';
          WHEN "110011" =>
            uut_h_0_0_i <= "000000000111111000001011100";
            uut_h_0_1_i <= "111111110101011001110001000";
            uut_h_0_2_i <= "111111110101011011000110101";
            uut_h_1_0_i <= "111111110011110000100111100";
            uut_h_1_1_i <= "000000001010100110000111011";
            uut_h_1_2_i <= "000000001100010001111001001";
            uut_coord_trans <= "111111101000";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111110101010100101100001" OR uut_h_0_1 /= "000000000001110100011110000010" OR uut_h_0_2 /= "000000000001111000111100000101" OR uut_h_1_0 /= "111111111110100110010011001010" OR uut_h_1_1 /= "111111111110000100000100101001" OR uut_h_1_2 /= "000000001111001110101011001100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "110000";
              state <= "111110";
            ELSE
              state <= "110100";
            END IF;
            uut_rst <= '0';
          WHEN "110100" =>
            uut_h_0_0_i <= "111111111000101011111011111";
            uut_h_0_1_i <= "111111111110010101001111100";
            uut_h_0_2_i <= "111111110101100100100101111";
            uut_h_1_0_i <= "000000001011110001011011001";
            uut_h_1_1_i <= "000000000110101101010101110";
            uut_h_1_2_i <= "111111110111110100111011101";
            uut_coord_trans <= "000000111101";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000001011100110000100100" OR uut_h_0_1 /= "000000000000101001001001001110" OR uut_h_0_2 /= "000000000010101000001101011101" OR uut_h_1_0 /= "000000000001100101011110101100" OR uut_h_1_1 /= "000000000001110000111101001000" OR uut_h_1_2 /= "000000111100001010100100100011" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "110001";
              state <= "111110";
            ELSE
              state <= "110101";
            END IF;
            uut_rst <= '0';
          WHEN "110101" =>
            uut_h_0_0_i <= "000000001011010011101101000";
            uut_h_0_1_i <= "111111110010100100011010100";
            uut_h_0_2_i <= "111111110110110111100001010";
            uut_h_1_0_i <= "111111111100101111010110000";
            uut_h_1_1_i <= "111111111011100010001111001";
            uut_h_1_2_i <= "000000001001010100000011001";
            uut_coord_trans <= "111110100001";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111110010010001111111011" OR uut_h_0_1 /= "000000000001111111001111100001" OR uut_h_0_2 /= "000001000010001100100101011100" OR uut_h_1_0 /= "111111111111111101001101110101" OR uut_h_1_1 /= "111111111110000001000111111101" OR uut_h_1_2 /= "000010011000100110111110100011" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "110010";
              state <= "111110";
            ELSE
              state <= "110110";
            END IF;
            uut_rst <= '0';
          WHEN "110110" =>
            uut_h_0_0_i <= "000000001001001001010001010";
            uut_h_0_1_i <= "000000001010101100000011100";
            uut_h_0_2_i <= "000000001101100111111010000";
            uut_h_1_0_i <= "000000001101100001011010001";
            uut_h_1_1_i <= "111111110100001101000000110";
            uut_h_1_2_i <= "000000001010101001011000101";
            uut_coord_trans <= "111111000110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000111111000001011100" OR uut_h_0_1 /= "111111111110101011001110001000" OR uut_h_0_2 /= "111111100010100110010011100101" OR uut_h_1_0 /= "111111111110011110000100111100" OR uut_h_1_1 /= "000000000001010100110000111011" OR uut_h_1_2 /= "111111100111000100010101011101" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "110011";
              state <= "111110";
            ELSE
              state <= "110111";
            END IF;
            uut_rst <= '0';
          WHEN "110111" =>
            uut_h_0_0_i <= "000000000000101101101100110";
            uut_h_0_1_i <= "000000001111110011100000111";
            uut_h_0_2_i <= "111111111111101100011011001";
            uut_h_1_0_i <= "111111111100101101110010011";
            uut_h_1_1_i <= "000000000011010101111110001";
            uut_h_1_2_i <= "111111111110000000111010100";
            uut_coord_trans <= "000000110000";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111111000101011111011111" OR uut_h_0_1 /= "111111111111110010101001111100" OR uut_h_0_2 /= "000001011101111100000101011000" OR uut_h_1_0 /= "000000000001011110001011011001" OR uut_h_1_1 /= "000000000000110101101010101110" OR uut_h_1_2 /= "111111110101100001010101001000" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "110100";
              state <= "111110";
            ELSE
              state <= "111000";
            END IF;
            uut_rst <= '0';
          WHEN "111000" =>
            uut_h_0_0_i <= "111111111110001011000100010";
            uut_h_0_1_i <= "000000001001100010010001100";
            uut_h_0_2_i <= "000000000001110100110111110";
            uut_h_1_0_i <= "111111110001101100100010110";
            uut_h_1_1_i <= "000000000100111110101000011";
            uut_h_1_2_i <= "000000000111000010001001110";
            uut_coord_trans <= "111111000111";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000001011010011101101000" OR uut_h_0_1 /= "111111111110010100100011010100" OR uut_h_0_2 /= "111110010011010000001000101100" OR uut_h_1_0 /= "111111111111100101111010110000" OR uut_h_1_1 /= "111111111111011100010001111001" OR uut_h_1_2 /= "111101110100010010111000110101" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "110101";
              state <= "111110";
            ELSE
              state <= "111001";
            END IF;
            uut_rst <= '0';
          WHEN "111001" =>
            uut_h_0_0_i <= "000000001001111100111110000";
            uut_h_0_1_i <= "000000001101100011011100010";
            uut_h_0_2_i <= "111111110101010111101011011";
            uut_h_1_0_i <= "111111110100011011111110101";
            uut_h_1_1_i <= "111111110000011010000111111";
            uut_h_1_2_i <= "000000000001010010011000000";
            uut_coord_trans <= "111110100011";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000001001001001010001010" OR uut_h_0_1 /= "000000000001010101100000011100" OR uut_h_0_2 /= "000000001111100110010010011110" OR uut_h_1_0 /= "000000000001101100001011010001" OR uut_h_1_1 /= "111111111110100001101000000110" OR uut_h_1_2 /= "111111001101100101011100100000" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "110110";
              state <= "111110";
            ELSE
              state <= "111010";
            END IF;
            uut_rst <= '0';
          WHEN "111010" =>
            uut_h_0_0_i <= "000000001101110111010000001";
            uut_h_0_1_i <= "000000000100100111010101010";
            uut_h_0_2_i <= "111111110001010001000110111";
            uut_h_1_0_i <= "000000001111000101110100011";
            uut_h_1_1_i <= "111111110010001011001001111";
            uut_h_1_2_i <= "111111111111000001001111110";
            uut_coord_trans <= "000001100010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000000000101101101100110" OR uut_h_0_1 /= "000000000001111110011100000111" OR uut_h_0_2 /= "111111111110011001111010100001" OR uut_h_1_0 /= "111111111111100101101110010011" OR uut_h_1_1 /= "000000000000011010101111110001" OR uut_h_1_2 /= "000000101111100100110101110100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "110111";
              state <= "111110";
            ELSE
              state <= "111011";
            END IF;
            uut_rst <= '0';
          WHEN "111011" =>
            IF uut_h_0_0 /= "111111111111110001011000100010" OR uut_h_0_1 /= "000000000001001100010010001100" OR uut_h_0_2 /= "111111100010101100001000011101" OR uut_h_1_0 /= "111111111110001101100100010110" OR uut_h_1_1 /= "000000000000100111110101000011" OR uut_h_1_2 /= "111110100110101010000100110111" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "111000";
              state <= "111110";
            ELSE
              state <= "111100";
            END IF;
            uut_rst <= '0';
          WHEN "111100" =>
            IF uut_h_0_0 /= "000000000001001111100111110000" OR uut_h_0_1 /= "000000000001101100011011100010" OR uut_h_0_2 /= "000000101010010011010110000000" OR uut_h_1_0 /= "111111111110100011011111110101" OR uut_h_1_1 /= "111111111110000011010000111111" OR uut_h_1_2 /= "111100000101010100110000110011" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "111001";
              state <= "111110";
            ELSE
              state <= "111101";
            END IF;
            uut_rst <= '0';
          WHEN "111101" =>
            IF uut_h_0_0 /= "000000000001101110111010000001" OR uut_h_0_1 /= "000000000000100100111010101010" OR uut_h_0_2 /= "111111101110111110110011111100" OR uut_h_1_0 /= "000000000001111000101110100011" OR uut_h_1_1 /= "111111111110010001011001001111" OR uut_h_1_2 /= "000001011010001000001100101100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "111010";
              state <= "111110";
            ELSE
              state <= "111110";
            END IF;
            uut_rst <= '0';
          WHEN OTHERS =>
            DONE <= '1';
            uut_rst <= '1';
        END CASE;
      END IF;
    END IF;
  END PROCESS;
END;
