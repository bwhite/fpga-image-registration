/home/brandyn/fpga-image-registration/modules/./fetch_stage/fetch_stage.vhd