/home/brandyn/fpga-image-registration/modules/./compose_h_matrix/compose_h_matrix.vhd