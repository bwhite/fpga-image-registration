LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
ENTITY affine_coord_transformT0_tb IS
PORT(
  CLK : IN STD_LOGIC;
  RST : IN STD_LOGIC;
  DONE : OUT STD_LOGIC;
  FAIL : OUT STD_LOGIC;
  FAIL_NUM : OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END affine_coord_transformT0_tb;
ARCHITECTURE behavior OF affine_coord_transformT0_tb IS
  COMPONENT affine_coord_transform
  PORT(
    CLK : IN STD_LOGIC;
    RST : IN STD_LOGIC;
    INPUT_VALID : IN STD_LOGIC;
    X_COORD : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    Y_COORD : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    H_0_0 : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    H_1_0 : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    H_0_1 : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    H_1_1 : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    H_0_2 : IN STD_LOGIC_VECTOR(21 DOWNTO 0);
    H_1_2 : IN STD_LOGIC_VECTOR(21 DOWNTO 0);
    XP_COORD : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
    YP_COORD : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
    OVERFLOW_X : OUT STD_LOGIC;
    OVERFLOW_Y : OUT STD_LOGIC;
    OUTPUT_VALID : OUT STD_LOGIC);
  END COMPONENT;
  SIGNAL uut_rst_wire, uut_rst : STD_LOGIC;
  SIGNAL state : STD_LOGIC_VECTOR(6 DOWNTO 0);
  -- UUT Input
  SIGNAL uut_input_valid : STD_LOGIC;
  SIGNAL uut_x_coord, uut_y_coord : STD_LOGIC_VECTOR(9 DOWNTO 0);
  SIGNAL uut_h_0_0, uut_h_1_0, uut_h_0_1, uut_h_1_1 : STD_LOGIC_VECTOR(17 DOWNTO 0);
  SIGNAL uut_h_0_2, uut_h_1_2 : STD_LOGIC_VECTOR(21 DOWNTO 0);
  -- UUT Output
  SIGNAL uut_overflow_x, uut_overflow_y, uut_output_valid : STD_LOGIC;
  SIGNAL uut_xp_coord, uut_yp_coord : STD_LOGIC_VECTOR(9 DOWNTO 0);
BEGIN
  uut_rst_wire <= RST OR uut_rst;
  uut :  affine_coord_transform PORT MAP (
    CLK => CLK,
    RST => uut_rst_wire,
    INPUT_VALID => uut_input_valid,
    X_COORD => uut_x_coord,
    Y_COORD => uut_y_coord,
    H_0_0 => uut_h_0_0,
    H_1_0 => uut_h_1_0,
    H_0_1 => uut_h_0_1,
    H_1_1 => uut_h_1_1,
    H_0_2 => uut_h_0_2,
    H_1_2 => uut_h_1_2,
    XP_COORD => uut_xp_coord,
    YP_COORD => uut_yp_coord,
    OVERFLOW_X => uut_overflow_x,
    OVERFLOW_Y => uut_overflow_y,
    OUTPUT_VALID => uut_output_valid
  );
  PROCESS (CLK) IS
  BEGIN
    IF CLK'event AND CLK='1' THEN
      IF RST='1' THEN
        DONE <= '0';
        FAIL <= '0';
        uut_rst <= '1';
        FAIL_NUM <= (OTHERS => '0');
        state <= (OTHERS => '0');
      ELSE
        CASE state IS
          WHEN "0000000" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0010110111";
            uut_y_coord <= "0100010001";
            uut_h_0_0 <= "000000100000000000";
            uut_h_1_0 <= "000000000000000000";
            uut_h_0_1 <= "000000000000000000";
            uut_h_1_1 <= "000000100000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            state <= "0000001";
            uut_rst <= '0';
          WHEN "0000001" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0000000110";
            uut_y_coord <= "0010100010";
            uut_h_0_0 <= "000000100000000000";
            uut_h_1_0 <= "000000000000000000";
            uut_h_0_1 <= "000000000000000000";
            uut_h_1_1 <= "000000100000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            state <= "0000010";
            uut_rst <= '0';
          WHEN "0000010" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0101001011";
            uut_y_coord <= "0101100111";
            uut_h_0_0 <= "000000100000000000";
            uut_h_1_0 <= "000000000000000000";
            uut_h_0_1 <= "000000000000000000";
            uut_h_1_1 <= "000000100000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            state <= "0000011";
            uut_rst <= '0';
          WHEN "0000011" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0000100110";
            uut_y_coord <= "0011010100";
            uut_h_0_0 <= "000000100000000000";
            uut_h_1_0 <= "000000000000000000";
            uut_h_0_1 <= "000000000000000000";
            uut_h_1_1 <= "000000100000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            state <= "0000100";
            uut_rst <= '0';
          WHEN "0000100" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0001111101";
            uut_y_coord <= "0110000000";
            uut_h_0_0 <= "000000100000000000";
            uut_h_1_0 <= "000000000000000000";
            uut_h_0_1 <= "000000000000000000";
            uut_h_1_1 <= "000000100000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            state <= "0000101";
            uut_rst <= '0';
          WHEN "0000101" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0100001000";
            uut_y_coord <= "0001000110";
            uut_h_0_0 <= "000000100000000000";
            uut_h_1_0 <= "000000000000000000";
            uut_h_0_1 <= "000000000000000000";
            uut_h_1_1 <= "000000100000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0010110111" OR uut_yp_coord /= "0100010001" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0000000";
              state <= "1011101";
            ELSE
              state <= "0000110";
            END IF;
            uut_rst <= '0';
          WHEN "0000110" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0110101101";
            uut_y_coord <= "0101010010";
            uut_h_0_0 <= "000000000000000000";
            uut_h_1_0 <= "000000100000000000";
            uut_h_0_1 <= "000000100000000000";
            uut_h_1_1 <= "000000000000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0000000110" OR uut_yp_coord /= "0010100010" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0000001";
              state <= "1011101";
            ELSE
              state <= "0000111";
            END IF;
            uut_rst <= '0';
          WHEN "0000111" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0001010000";
            uut_y_coord <= "0100101011";
            uut_h_0_0 <= "000000000000000000";
            uut_h_1_0 <= "000000100000000000";
            uut_h_0_1 <= "000000100000000000";
            uut_h_1_1 <= "000000000000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0101001011" OR uut_yp_coord /= "0101100111" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0000010";
              state <= "1011101";
            ELSE
              state <= "0001000";
            END IF;
            uut_rst <= '0';
          WHEN "0001000" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0011000001";
            uut_y_coord <= "0100101010";
            uut_h_0_0 <= "000000000000000000";
            uut_h_1_0 <= "000000100000000000";
            uut_h_0_1 <= "000000100000000000";
            uut_h_1_1 <= "000000000000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0000100110" OR uut_yp_coord /= "0011010100" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0000011";
              state <= "1011101";
            ELSE
              state <= "0001001";
            END IF;
            uut_rst <= '0';
          WHEN "0001001" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0011111111";
            uut_y_coord <= "0110010000";
            uut_h_0_0 <= "000000000000000000";
            uut_h_1_0 <= "000000100000000000";
            uut_h_0_1 <= "000000100000000000";
            uut_h_1_1 <= "000000000000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0001111101" OR uut_yp_coord /= "0110000000" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0000100";
              state <= "1011101";
            ELSE
              state <= "0001010";
            END IF;
            uut_rst <= '0';
          WHEN "0001010" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0011001100";
            uut_y_coord <= "0011001110";
            uut_h_0_0 <= "000000000000000000";
            uut_h_1_0 <= "000000100000000000";
            uut_h_0_1 <= "000000100000000000";
            uut_h_1_1 <= "000000000000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0100001000" OR uut_yp_coord /= "0001000110" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0000101";
              state <= "1011101";
            ELSE
              state <= "0001011";
            END IF;
            uut_rst <= '0';
          WHEN "0001011" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0001110011";
            uut_y_coord <= "0101101111";
            uut_h_0_0 <= "000000000000000000";
            uut_h_1_0 <= "000000100000000000";
            uut_h_0_1 <= "000000100000000000";
            uut_h_1_1 <= "000000000000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0101010010" OR uut_yp_coord /= "0110101101" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0000110";
              state <= "1011101";
            ELSE
              state <= "0001100";
            END IF;
            uut_rst <= '0';
          WHEN "0001100" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0110001011";
            uut_y_coord <= "0001010100";
            uut_h_0_0 <= "000000000000000000";
            uut_h_1_0 <= "000000100000000000";
            uut_h_0_1 <= "000000100000000000";
            uut_h_1_1 <= "000000000000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0100101011" OR uut_yp_coord /= "0001010000" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0000111";
              state <= "1011101";
            ELSE
              state <= "0001101";
            END IF;
            uut_rst <= '0';
          WHEN "0001101" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0101000110";
            uut_y_coord <= "0000010010";
            uut_h_0_0 <= "000000000000000000";
            uut_h_1_0 <= "000000100000000000";
            uut_h_0_1 <= "000000100000000000";
            uut_h_1_1 <= "000000000000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0100101010" OR uut_yp_coord /= "0011000001" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0001000";
              state <= "1011101";
            ELSE
              state <= "0001110";
            END IF;
            uut_rst <= '0';
          WHEN "0001110" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0001010111";
            uut_y_coord <= "0001111011";
            uut_h_0_0 <= "000000000000000000";
            uut_h_1_0 <= "000000100000000000";
            uut_h_0_1 <= "000000100000000000";
            uut_h_1_1 <= "000000000000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0110010000" OR uut_yp_coord /= "0011111111" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0001001";
              state <= "1011101";
            ELSE
              state <= "0001111";
            END IF;
            uut_rst <= '0';
          WHEN "0001111" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0011010011";
            uut_y_coord <= "0001111100";
            uut_h_0_0 <= "000000000000000000";
            uut_h_1_0 <= "000000100000000000";
            uut_h_0_1 <= "000000100000000000";
            uut_h_1_1 <= "000000000000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0011001110" OR uut_yp_coord /= "0011001100" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0001010";
              state <= "1011101";
            ELSE
              state <= "0010000";
            END IF;
            uut_rst <= '0';
          WHEN "0010000" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0010111100";
            uut_y_coord <= "0110001000";
            uut_h_0_0 <= "000000000000000000";
            uut_h_1_0 <= "000000100000000000";
            uut_h_0_1 <= "000000100000000000";
            uut_h_1_1 <= "000000000000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0101101111" OR uut_yp_coord /= "0001110011" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0001011";
              state <= "1011101";
            ELSE
              state <= "0010001";
            END IF;
            uut_rst <= '0';
          WHEN "0010001" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0000011101";
            uut_y_coord <= "0110100000";
            uut_h_0_0 <= "000000000000000000";
            uut_h_1_0 <= "000000100000000000";
            uut_h_0_1 <= "000000100000000000";
            uut_h_1_1 <= "000000000000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0001010100" OR uut_yp_coord /= "0110001011" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0001100";
              state <= "1011101";
            ELSE
              state <= "0010010";
            END IF;
            uut_rst <= '0';
          WHEN "0010010" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0000001100";
            uut_y_coord <= "0011001010";
            uut_h_0_0 <= "000000000000000000";
            uut_h_1_0 <= "000000100000000000";
            uut_h_0_1 <= "000000100000000000";
            uut_h_1_1 <= "000000000000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0000010010" OR uut_yp_coord /= "0101000110" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0001101";
              state <= "1011101";
            ELSE
              state <= "0010011";
            END IF;
            uut_rst <= '0';
          WHEN "0010011" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0001111111";
            uut_y_coord <= "0110111100";
            uut_h_0_0 <= "000000000000000000";
            uut_h_1_0 <= "000000100000000000";
            uut_h_0_1 <= "000000100000000000";
            uut_h_1_1 <= "000000000000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0001111011" OR uut_yp_coord /= "0001010111" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0001110";
              state <= "1011101";
            ELSE
              state <= "0010100";
            END IF;
            uut_rst <= '0';
          WHEN "0010100" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0100111101";
            uut_y_coord <= "0010111000";
            uut_h_0_0 <= "000000000000000000";
            uut_h_1_0 <= "000000100000000000";
            uut_h_0_1 <= "000000100000000000";
            uut_h_1_1 <= "000000000000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0001111100" OR uut_yp_coord /= "0011010011" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0001111";
              state <= "1011101";
            ELSE
              state <= "0010101";
            END IF;
            uut_rst <= '0';
          WHEN "0010101" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0100010100";
            uut_y_coord <= "0011111110";
            uut_h_0_0 <= "000000000000000000";
            uut_h_1_0 <= "000000100000000000";
            uut_h_0_1 <= "000000100000000000";
            uut_h_1_1 <= "000000000000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0110001000" OR uut_yp_coord /= "0010111100" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0010000";
              state <= "1011101";
            ELSE
              state <= "0010110";
            END IF;
            uut_rst <= '0';
          WHEN "0010110" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0000101010";
            uut_y_coord <= "0110000001";
            uut_h_0_0 <= "000000000000000000";
            uut_h_1_0 <= "000000100000000000";
            uut_h_0_1 <= "000000100000000000";
            uut_h_1_1 <= "000000000000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0110100000" OR uut_yp_coord /= "0000011101" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0010001";
              state <= "1011101";
            ELSE
              state <= "0010111";
            END IF;
            uut_rst <= '0';
          WHEN "0010111" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0110110000";
            uut_y_coord <= "0100101100";
            uut_h_0_0 <= "000000000000000000";
            uut_h_1_0 <= "000000100000000000";
            uut_h_0_1 <= "000000100000000000";
            uut_h_1_1 <= "000000000000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0011001010" OR uut_yp_coord /= "0000001100" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0010010";
              state <= "1011101";
            ELSE
              state <= "0011000";
            END IF;
            uut_rst <= '0';
          WHEN "0011000" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0011000101";
            uut_y_coord <= "0111011000";
            uut_h_0_0 <= "000000000000000000";
            uut_h_1_0 <= "000000100000000000";
            uut_h_0_1 <= "000000100000000000";
            uut_h_1_1 <= "000000000000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0110111100" OR uut_yp_coord /= "0001111111" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0010011";
              state <= "1011101";
            ELSE
              state <= "0011001";
            END IF;
            uut_rst <= '0';
          WHEN "0011001" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0101000110";
            uut_y_coord <= "0011111101";
            uut_h_0_0 <= "000000000000000000";
            uut_h_1_0 <= "000000100000000000";
            uut_h_0_1 <= "000000100000000000";
            uut_h_1_1 <= "000000000000000000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0010111000" OR uut_yp_coord /= "0100111101" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0010100";
              state <= "1011101";
            ELSE
              state <= "0011010";
            END IF;
            uut_rst <= '0';
          WHEN "0011010" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0001110010";
            uut_y_coord <= "0100010101";
            uut_h_0_0 <= "000000101001100110";
            uut_h_1_0 <= "000000101100110011";
            uut_h_0_1 <= "000000011100110011";
            uut_h_1_1 <= "000000100011001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0011111110" OR uut_yp_coord /= "0100010100" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0010101";
              state <= "1011101";
            ELSE
              state <= "0011011";
            END IF;
            uut_rst <= '0';
          WHEN "0011011" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0010111011";
            uut_y_coord <= "0010101101";
            uut_h_0_0 <= "000000101001100110";
            uut_h_1_0 <= "000000101100110011";
            uut_h_0_1 <= "000000011100110011";
            uut_h_1_1 <= "000000100011001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0110000001" OR uut_yp_coord /= "0000101010" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0010110";
              state <= "1011101";
            ELSE
              state <= "0011100";
            END IF;
            uut_rst <= '0';
          WHEN "0011100" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0011101101";
            uut_y_coord <= "0101010011";
            uut_h_0_0 <= "000000101001100110";
            uut_h_1_0 <= "000000101100110011";
            uut_h_0_1 <= "000000011100110011";
            uut_h_1_1 <= "000000100011001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0100101100" OR uut_yp_coord /= "0110110000" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0010111";
              state <= "1011101";
            ELSE
              state <= "0011101";
            END IF;
            uut_rst <= '0';
          WHEN "0011101" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0001000100";
            uut_y_coord <= "0010000000";
            uut_h_0_0 <= "000000101001100110";
            uut_h_1_0 <= "000000101100110011";
            uut_h_0_1 <= "000000011100110011";
            uut_h_1_1 <= "000000100011001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0111011000" OR uut_yp_coord /= "0011000101" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0011000";
              state <= "1011101";
            ELSE
              state <= "0011110";
            END IF;
            uut_rst <= '0';
          WHEN "0011110" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0011111011";
            uut_y_coord <= "0001111111";
            uut_h_0_0 <= "000000101001100110";
            uut_h_1_0 <= "000000101100110011";
            uut_h_0_1 <= "000000011100110011";
            uut_h_1_1 <= "000000100011001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0011111101" OR uut_yp_coord /= "0101000110" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0011001";
              state <= "1011101";
            ELSE
              state <= "0011111";
            END IF;
            uut_rst <= '0';
          WHEN "0011111" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0000000011";
            uut_y_coord <= "0101000110";
            uut_h_0_0 <= "000000101001100110";
            uut_h_1_0 <= "000000101100110011";
            uut_h_0_1 <= "000000011100110011";
            uut_h_1_1 <= "000000100011001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0110001101" OR uut_yp_coord /= "0111010000" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0011010";
              state <= "1011101";
            ELSE
              state <= "0100000";
            END IF;
            uut_rst <= '0';
          WHEN "0100000" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0110011011";
            uut_y_coord <= "0011000001";
            uut_h_0_0 <= "000000101001100110";
            uut_h_1_0 <= "000000101100110011";
            uut_h_0_1 <= "000000011100110011";
            uut_h_1_1 <= "000000100011001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0110001110" OR uut_yp_coord /= "0111000100" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0011011";
              state <= "1011101";
            ELSE
              state <= "0100001";
            END IF;
            uut_rst <= '0';
          WHEN "0100001" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0110110010";
            uut_y_coord <= "0000001111";
            uut_h_0_0 <= "000000101001100110";
            uut_h_1_0 <= "000000101100110011";
            uut_h_0_1 <= "000000011100110011";
            uut_h_1_1 <= "000000100011001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "1001100101" OR uut_yp_coord /= "1011000000" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0011100";
              state <= "1011101";
            ELSE
              state <= "0100010";
            END IF;
            uut_rst <= '0';
          WHEN "0100010" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0000010111";
            uut_y_coord <= "0100001001";
            uut_h_0_0 <= "000000101001100110";
            uut_h_1_0 <= "000000101100110011";
            uut_h_0_1 <= "000000011100110011";
            uut_h_1_1 <= "000000100011001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0011001011" OR uut_yp_coord /= "0011101011" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0011101";
              state <= "1011101";
            ELSE
              state <= "0100011";
            END IF;
            uut_rst <= '0';
          WHEN "0100011" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0001010100";
            uut_y_coord <= "0010101100";
            uut_h_0_0 <= "000000101001100110";
            uut_h_1_0 <= "000000101100110011";
            uut_h_0_1 <= "000000011100110011";
            uut_h_1_1 <= "000000100011001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0110111000" OR uut_yp_coord /= "0111101011" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0011110";
              state <= "1011101";
            ELSE
              state <= "0100100";
            END IF;
            uut_rst <= '0';
          WHEN "0100100" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0011110000";
            uut_y_coord <= "0101101101";
            uut_h_0_0 <= "000000101001100110";
            uut_h_1_0 <= "000000101100110011";
            uut_h_0_1 <= "000000011100110011";
            uut_h_1_1 <= "000000100011001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0100101001" OR uut_yp_coord /= "0101101010" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0011111";
              state <= "1011101";
            ELSE
              state <= "0100101";
            END IF;
            uut_rst <= '0';
          WHEN "0100101" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0001000110";
            uut_y_coord <= "0001011111";
            uut_h_0_0 <= "000000101001100110";
            uut_h_1_0 <= "000000101100110011";
            uut_h_0_1 <= "000000011100110011";
            uut_h_1_1 <= "000000100011001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "1011000011" OR uut_yp_coord /= "1100010011" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0100000";
              state <= "1011101";
            ELSE
              state <= "0100110";
            END IF;
            uut_rst <= '0';
          WHEN "0100110" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0110110011";
            uut_y_coord <= "0010111100";
            uut_h_0_0 <= "000000101001100110";
            uut_h_1_0 <= "000000101100110011";
            uut_h_0_1 <= "000000011100110011";
            uut_h_1_1 <= "000000100011001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "1001000001" OR uut_yp_coord /= "1001110000" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0100001";
              state <= "1011101";
            ELSE
              state <= "0100111";
            END IF;
            uut_rst <= '0';
          WHEN "0100111" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0101011001";
            uut_y_coord <= "0100111000";
            uut_h_0_0 <= "000000101001100110";
            uut_h_1_0 <= "000000101100110011";
            uut_h_0_1 <= "000000011100110011";
            uut_h_1_1 <= "000000100011001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0100001100" OR uut_yp_coord /= "0101000011" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0100010";
              state <= "1011101";
            ELSE
              state <= "0101000";
            END IF;
            uut_rst <= '0';
          WHEN "0101000" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0111001101";
            uut_y_coord <= "0001011001";
            uut_h_0_0 <= "000000101001100110";
            uut_h_1_0 <= "000000101100110011";
            uut_h_0_1 <= "000000011100110011";
            uut_h_1_1 <= "000000100011001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0100000111" OR uut_yp_coord /= "0100110010" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0100011";
              state <= "1011101";
            ELSE
              state <= "0101001";
            END IF;
            uut_rst <= '0';
          WHEN "0101001" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0000111110";
            uut_y_coord <= "0011010000";
            uut_h_0_0 <= "000000101001100110";
            uut_h_1_0 <= "000000101100110011";
            uut_h_0_1 <= "000000011100110011";
            uut_h_1_1 <= "000000100011001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "1010000000" OR uut_yp_coord /= "1011100001" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0100100";
              state <= "1011101";
            ELSE
              state <= "0101010";
            END IF;
            uut_rst <= '0';
          WHEN "0101010" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0000011101";
            uut_y_coord <= "0011101110";
            uut_h_0_0 <= "000000101001100110";
            uut_h_1_0 <= "000000101100110011";
            uut_h_0_1 <= "000000011100110011";
            uut_h_1_1 <= "000000100011001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0010110000" OR uut_yp_coord /= "0011001010" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0100101";
              state <= "1011101";
            ELSE
              state <= "0101011";
            END IF;
            uut_rst <= '0';
          WHEN "0101011" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0001110001";
            uut_y_coord <= "0111001011";
            uut_h_0_0 <= "000000101001100110";
            uut_h_1_0 <= "000000101100110011";
            uut_h_0_1 <= "000000011100110011";
            uut_h_1_1 <= "000000100011001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "1011011110" OR uut_yp_coord /= "1100101111" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0100110";
              state <= "1011101";
            ELSE
              state <= "0101100";
            END IF;
            uut_rst <= '0';
          WHEN "0101100" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0101011100";
            uut_y_coord <= "0001101110";
            uut_h_0_0 <= "000000101001100110";
            uut_h_1_0 <= "000000101100110011";
            uut_h_0_1 <= "000000011100110011";
            uut_h_1_1 <= "000000100011001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "1011011001" OR uut_yp_coord /= "1100111010" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0100111";
              state <= "1011101";
            ELSE
              state <= "0101101";
            END IF;
            uut_rst <= '0';
          WHEN "0101101" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0101011100";
            uut_y_coord <= "0100001011";
            uut_h_0_0 <= "000000101001100110";
            uut_h_1_0 <= "000000101100110011";
            uut_h_0_1 <= "000000011100110011";
            uut_h_1_1 <= "000000100011001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "1010100111" OR uut_yp_coord /= "1011100111" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0101000";
              state <= "1011101";
            ELSE
              state <= "0101110";
            END IF;
            uut_rst <= '0';
          WHEN "0101110" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0101010100";
            uut_y_coord <= "0010010101";
            uut_h_0_0 <= "000000000111000001";
            uut_h_1_0 <= "000000010001010001";
            uut_h_0_1 <= "000000100001100100";
            uut_h_1_1 <= "000000111110001111";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0100001011" OR uut_yp_coord /= "0100111011" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0101001";
              state <= "1011101";
            ELSE
              state <= "0101111";
            END IF;
            uut_rst <= '0';
          WHEN "0101111" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0110001101";
            uut_y_coord <= "0001011011";
            uut_h_0_0 <= "000000111100101011";
            uut_h_1_0 <= "000000000011111001";
            uut_h_0_1 <= "000000100101011010";
            uut_h_1_1 <= "000000010010001111";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0011111011" OR uut_yp_coord /= "0100101110" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0101010";
              state <= "1011101";
            ELSE
              state <= "0110000";
            END IF;
            uut_rst <= '0';
          WHEN "0110000" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0110110011";
            uut_y_coord <= "0100001001";
            uut_h_0_0 <= "000000100100100010";
            uut_h_1_0 <= "000000001010110111";
            uut_h_0_1 <= "000000001001011100";
            uut_h_1_1 <= "000000011110011110";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "1000101111" OR uut_yp_coord /= "1010010110" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0101011";
              state <= "1011101";
            ELSE
              state <= "0110001";
            END IF;
            uut_rst <= '0';
          WHEN "0110001" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0111010011";
            uut_y_coord <= "0000100100";
            uut_h_0_0 <= "000000101101100010";
            uut_h_1_0 <= "000000110111110001";
            uut_h_0_1 <= "000000010101000010";
            uut_h_1_1 <= "000000101001100110";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "1000100111" OR uut_yp_coord /= "1001100000" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0101100";
              state <= "1011101";
            ELSE
              state <= "0110010";
            END IF;
            uut_rst <= '0';
          WHEN "0110010" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0101011101";
            uut_y_coord <= "0011101111";
            uut_h_0_0 <= "000000001100100001";
            uut_h_1_0 <= "000000111111100000";
            uut_h_0_1 <= "000000110011010110";
            uut_h_1_1 <= "000000011011001001";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "1010110100" OR uut_yp_coord /= "1100001100" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0101101";
              state <= "1011101";
            ELSE
              state <= "0110011";
            END IF;
            uut_rst <= '0';
          WHEN "0110011" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0001011000";
            uut_y_coord <= "0011101111";
            uut_h_0_0 <= "000000000010100000";
            uut_h_1_0 <= "000000111100100100";
            uut_h_0_1 <= "000000110000111000";
            uut_h_1_1 <= "000000100011110000";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0011100110" OR uut_yp_coord /= "0111011001" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0101110";
              state <= "1011101";
            ELSE
              state <= "0110100";
            END IF;
            uut_rst <= '0';
          WHEN "0110100" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0101101011";
            uut_y_coord <= "0111011101";
            uut_h_0_0 <= "000000001110110101";
            uut_h_1_0 <= "000000011001010111";
            uut_h_0_1 <= "000000101101000111";
            uut_h_1_1 <= "000000100011101111";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "1101011011" OR uut_yp_coord /= "0001100100" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0101111";
              state <= "1011101";
            ELSE
              state <= "0110101";
            END IF;
            uut_rst <= '0';
          WHEN "0110101" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0101010101";
            uut_y_coord <= "0000001000";
            uut_h_0_0 <= "000000111001101011";
            uut_h_1_0 <= "000000100010100110";
            uut_h_0_1 <= "000000011011101001";
            uut_h_1_1 <= "000000100010101110";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "1000111110" OR uut_yp_coord /= "0110001111" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0110000";
              state <= "1011101";
            ELSE
              state <= "0110110";
            END IF;
            uut_rst <= '0';
          WHEN "0110110" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0011100010";
            uut_y_coord <= "0011000001";
            uut_h_0_0 <= "000000001100101011";
            uut_h_1_0 <= "000000001100011111";
            uut_h_0_1 <= "000000010100111010";
            uut_h_1_1 <= "000000111000010101";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "1010110000" OR uut_yp_coord /= "1101011100" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0110001";
              state <= "1011101";
            ELSE
              state <= "0110111";
            END IF;
            uut_rst <= '0';
          WHEN "0110111" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0010100000";
            uut_y_coord <= "0100011110";
            uut_h_0_0 <= "000000011101110000";
            uut_h_1_0 <= "000000110100000110";
            uut_h_0_1 <= "000000111001100000";
            uut_h_1_1 <= "000000011011011110";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "1000000111" OR uut_yp_coord /= "1101111111" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0110010";
              state <= "1011101";
            ELSE
              state <= "0111000";
            END IF;
            uut_rst <= '0';
          WHEN "0111000" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0000000100";
            uut_y_coord <= "0110110111";
            uut_h_0_0 <= "000000000100100011";
            uut_h_1_0 <= "000000001011101001";
            uut_h_0_1 <= "000000000101111100";
            uut_h_1_1 <= "000000011101101010";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0101110011" OR uut_yp_coord /= "0110110001" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0110011";
              state <= "1011101";
            ELSE
              state <= "0111001";
            END IF;
            uut_rst <= '0';
          WHEN "0111001" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0000010111";
            uut_y_coord <= "0000010111";
            uut_h_0_0 <= "000000010110101010";
            uut_h_1_0 <= "000000110001111100";
            uut_h_0_1 <= "000000011011111100";
            uut_h_1_1 <= "000000011011111100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "1101001000" OR uut_yp_coord /= "1100110100" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0110100";
              state <= "1011101";
            ELSE
              state <= "0111010";
            END IF;
            uut_rst <= '0';
          WHEN "0111010" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0011011101";
            uut_y_coord <= "0100110010";
            uut_h_0_0 <= "000000001110011110";
            uut_h_1_0 <= "000000100010010110";
            uut_h_0_1 <= "000000110000110001";
            uut_h_1_1 <= "000000010110001111";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "1001101101" OR uut_yp_coord /= "0101111001" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0110101";
              state <= "1011101";
            ELSE
              state <= "0111011";
            END IF;
            uut_rst <= '0';
          WHEN "0111011" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0000111011";
            uut_y_coord <= "0011100001";
            uut_h_0_0 <= "000000010111100111";
            uut_h_1_0 <= "000000001101010101";
            uut_h_0_1 <= "000000011100001110";
            uut_h_1_1 <= "000000111101001100";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0011010111" OR uut_yp_coord /= "0110101011" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0110110";
              state <= "1011101";
            ELSE
              state <= "0111100";
            END IF;
            uut_rst <= '0';
          WHEN "0111100" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0010100110";
            uut_y_coord <= "0011001000";
            uut_h_0_0 <= "000000100111000110";
            uut_h_1_0 <= "000000111001100110";
            uut_h_0_1 <= "000000001100011000";
            uut_h_1_1 <= "000000110000010010";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "1010010110" OR uut_yp_coord /= "0111111001" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0110111";
              state <= "1011101";
            ELSE
              state <= "0111101";
            END IF;
            uut_rst <= '0';
          WHEN "0111101" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0011011011";
            uut_y_coord <= "0100101000";
            uut_h_0_0 <= "000000110000010101";
            uut_h_1_0 <= "000000101111100000";
            uut_h_0_1 <= "000000110101001100";
            uut_h_1_1 <= "000000001010000001";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0001010010" OR uut_yp_coord /= "0110011000" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0111000";
              state <= "1011101";
            ELSE
              state <= "0111110";
            END IF;
            uut_rst <= '0';
          WHEN "0111110" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0001000101";
            uut_y_coord <= "0100100010";
            uut_h_0_0 <= "000000011010000110";
            uut_h_1_0 <= "000000000010010101";
            uut_h_0_1 <= "000000101111110000";
            uut_h_1_1 <= "000000001001111010";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0000100100" OR uut_yp_coord /= "0000110111" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0111001";
              state <= "1011101";
            ELSE
              state <= "0111111";
            END IF;
            uut_rst <= '0';
          WHEN "0111111" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0101100011";
            uut_y_coord <= "0101001100";
            uut_h_0_0 <= "000000000110000011";
            uut_h_1_0 <= "000000010100101011";
            uut_h_0_1 <= "000000110001010000";
            uut_h_1_1 <= "000000001110111110";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "1000110110" OR uut_yp_coord /= "0111000001" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0111010";
              state <= "1011101";
            ELSE
              state <= "1000000";
            END IF;
            uut_rst <= '0';
          WHEN "1000000" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0011011011";
            uut_y_coord <= "0010111000";
            uut_h_0_0 <= "000000100011101001";
            uut_h_1_0 <= "000000010000110101";
            uut_h_0_1 <= "000000101011100011";
            uut_h_1_1 <= "000000001110111101";
            uut_h_0_2 <= "0000000000000000000000";
            uut_h_1_2 <= "0000000000000000000000";
            IF uut_xp_coord /= "0011110001" OR uut_yp_coord /= "0111000110" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0111011";
              state <= "1011101";
            ELSE
              state <= "1000001";
            END IF;
            uut_rst <= '0';
          WHEN "1000001" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0100000011";
            uut_y_coord <= "0001100011";
            uut_h_0_0 <= "000000010011010000";
            uut_h_1_0 <= "000000011011011011";
            uut_h_0_1 <= "000000011111100111";
            uut_h_1_1 <= "000000011101101111";
            uut_h_0_2 <= "0001100010010010001001";
            uut_h_1_2 <= "0000000000000101001111";
            IF uut_xp_coord /= "0100011000" OR uut_yp_coord /= "1001011000" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0111100";
              state <= "1011101";
            ELSE
              state <= "1000010";
            END IF;
            uut_rst <= '0';
          WHEN "1000010" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0100101010";
            uut_y_coord <= "0101111110";
            uut_h_0_0 <= "000000010001101011";
            uut_h_1_0 <= "000000011110101001";
            uut_h_0_1 <= "000000011100100100";
            uut_h_1_1 <= "000000001011011010";
            uut_h_0_2 <= "0010000011001000101110";
            uut_h_1_2 <= "0001010011001101000010";
            IF uut_xp_coord /= "1100110110" OR uut_yp_coord /= "0110100001" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0111101";
              state <= "1011101";
            ELSE
              state <= "1000011";
            END IF;
            uut_rst <= '0';
          WHEN "1000011" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0010001001";
            uut_y_coord <= "0110111101";
            uut_h_0_0 <= "000000010111110101";
            uut_h_1_0 <= "000000011100100011";
            uut_h_0_1 <= "000000000111110000";
            uut_h_1_1 <= "000000000100001001";
            uut_h_0_2 <= "0000110110000001000010";
            uut_h_1_2 <= "0001010100000000001101";
            IF uut_xp_coord /= "0111101000" OR uut_yp_coord /= "0001011110" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0111110";
              state <= "1011101";
            ELSE
              state <= "1000100";
            END IF;
            uut_rst <= '0';
          WHEN "1000100" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0101000111";
            uut_y_coord <= "0111001101";
            uut_h_0_0 <= "000000000001100000";
            uut_h_1_0 <= "000000000110110101";
            uut_h_0_1 <= "000000001100101110";
            uut_h_1_1 <= "000000001010101011";
            uut_h_0_2 <= "0000110111000110101100";
            uut_h_1_2 <= "0011100000101010110011";
            IF uut_xp_coord /= "1001000010" OR uut_yp_coord /= "0110000000" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0111111";
              state <= "1011101";
            ELSE
              state <= "1000101";
            END IF;
            uut_rst <= '0';
          WHEN "1000101" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0100011000";
            uut_y_coord <= "0110001110";
            uut_h_0_0 <= "000000011010011100";
            uut_h_1_0 <= "000000010010010110";
            uut_h_0_1 <= "000000011001010111";
            uut_h_1_1 <= "000000001010100001";
            uut_h_0_2 <= "0000110101101000011000";
            uut_h_1_2 <= "0001001010111110010000";
            IF uut_xp_coord /= "0111101110" OR uut_yp_coord /= "0011001001" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1000000";
              state <= "1011101";
            ELSE
              state <= "1000110";
            END IF;
            uut_rst <= '0';
          WHEN "1000110" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0110001010";
            uut_y_coord <= "0110010011";
            uut_h_0_0 <= "000000000111111101";
            uut_h_1_0 <= "000000001111001110";
            uut_h_0_1 <= "000000001100110001";
            uut_h_1_1 <= "000000010011001011";
            uut_h_0_2 <= "0011000000001000000001";
            uut_h_1_2 <= "0000011001001101110110";
            IF uut_xp_coord /= "0111000010" OR uut_yp_coord /= "0100111010" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1000001";
              state <= "1011101";
            ELSE
              state <= "1000111";
            END IF;
            uut_rst <= '0';
          WHEN "1000111" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0111001110";
            uut_y_coord <= "0000101001";
            uut_h_0_0 <= "000000011110100110";
            uut_h_1_0 <= "000000010010010101";
            uut_h_0_1 <= "000000011011001100";
            uut_h_1_1 <= "000000001000110101";
            uut_h_0_2 <= "0010010101010110111001";
            uut_h_1_2 <= "0010001101001101001111";
            IF uut_xp_coord /= "1011111111" OR uut_yp_coord /= "1001001011" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1000010";
              state <= "1011101";
            ELSE
              state <= "1001000";
            END IF;
            uut_rst <= '0';
          WHEN "1001000" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0011100111";
            uut_y_coord <= "0010100010";
            uut_h_0_0 <= "000000010011110101";
            uut_h_1_0 <= "000000001000010101";
            uut_h_0_1 <= "000000001110010000";
            uut_h_1_1 <= "000000011011000000";
            uut_h_0_2 <= "0000101111000101101101";
            uut_h_1_2 <= "0001001000111011001010";
            IF uut_xp_coord /= "0100111101" OR uut_yp_coord /= "0101011011" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1000011";
              state <= "1011101";
            ELSE
              state <= "1001001";
            END IF;
            uut_rst <= '0';
          WHEN "1001001" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0111000000";
            uut_y_coord <= "0101011001";
            uut_h_0_0 <= "000000010100100110";
            uut_h_1_0 <= "000000011011100001";
            uut_h_0_1 <= "000000001100110111";
            uut_h_1_1 <= "000000010100001110";
            uut_h_0_2 <= "0011101100011101001111";
            uut_h_1_2 <= "0010000110010001100100";
            IF uut_xp_coord /= "0100110100" OR uut_yp_coord /= "1010100000" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1000100";
              state <= "1011101";
            ELSE
              state <= "1001010";
            END IF;
            uut_rst <= '0';
          WHEN "1001010" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0100010000";
            uut_y_coord <= "0111001101";
            uut_h_0_0 <= "000000011100110101";
            uut_h_1_0 <= "000000011111110110";
            uut_h_0_1 <= "000000010100111001";
            uut_h_1_1 <= "000000000011011110";
            uut_h_0_2 <= "0000001000101010101101";
            uut_h_1_2 <= "0010010100010101111000";
            IF uut_xp_coord /= "1010001101" OR uut_yp_coord /= "0110111001" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1000101";
              state <= "1011101";
            ELSE
              state <= "1001011";
            END IF;
            uut_rst <= '0';
          WHEN "1001011" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0010010101";
            uut_y_coord <= "0001101101";
            uut_h_0_0 <= "000000010000101000";
            uut_h_1_0 <= "000000000001111000";
            uut_h_0_1 <= "000000011100011110";
            uut_h_1_1 <= "000000001010100100";
            uut_h_0_2 <= "0000110111001000001101";
            uut_h_1_2 <= "0000011011010110010000";
            IF uut_xp_coord /= "1010000010" OR uut_yp_coord /= "0111011111" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1000110";
              state <= "1011101";
            ELSE
              state <= "1001100";
            END IF;
            uut_rst <= '0';
          WHEN "1001100" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0010011100";
            uut_y_coord <= "0100101110";
            uut_h_0_0 <= "000000011001000100";
            uut_h_1_0 <= "000000000011101001";
            uut_h_0_1 <= "000000011111010100";
            uut_h_1_1 <= "000000011011001001";
            uut_h_0_2 <= "0000001100001001111011";
            uut_h_1_2 <= "0001101111111000110111";
            IF uut_xp_coord /= "1100000111" OR uut_yp_coord /= "1000101110" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1000111";
              state <= "1011101";
            ELSE
              state <= "1001101";
            END IF;
            uut_rst <= '0';
          WHEN "1001101" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0110100010";
            uut_y_coord <= "0000011001";
            uut_h_0_0 <= "000000000011011101";
            uut_h_1_0 <= "000000001110101101";
            uut_h_0_1 <= "000000001110011011";
            uut_h_1_1 <= "000000010001101000";
            uut_h_0_2 <= "0011000001010011000000";
            uut_h_1_2 <= "0010101000001101000011";
            IF uut_xp_coord /= "0100110101" OR uut_yp_coord /= "0101010110" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1001000";
              state <= "1011101";
            ELSE
              state <= "1001110";
            END IF;
            uut_rst <= '0';
          WHEN "1001110" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0111000100";
            uut_y_coord <= "0000001000";
            uut_h_0_0 <= "000000010000001101";
            uut_h_1_0 <= "000000000110011001";
            uut_h_0_1 <= "000000001101101010";
            uut_h_1_1 <= "000000000101011001";
            uut_h_0_2 <= "0010110100011010000001";
            uut_h_1_2 <= "0001011000011001110111";
            IF uut_xp_coord /= "1110000011" OR uut_yp_coord /= "1101100111" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1001001";
              state <= "1011101";
            ELSE
              state <= "1001111";
            END IF;
            uut_rst <= '0';
          WHEN "1001111" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0100111000";
            uut_y_coord <= "0110011111";
            uut_h_0_0 <= "000000001001011010";
            uut_h_1_0 <= "000000000101110000";
            uut_h_0_1 <= "000000011101101001";
            uut_h_1_1 <= "000000000010001011";
            uut_h_0_2 <= "0010001011011101100101";
            uut_h_1_2 <= "0010011000111010101001";
            IF uut_xp_coord /= "1000110011" OR uut_yp_coord /= "1001101001" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1001010";
              state <= "1011101";
            ELSE
              state <= "1010000";
            END IF;
            uut_rst <= '0';
          WHEN "1010000" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0010100101";
            uut_y_coord <= "0111000110";
            uut_h_0_0 <= "000000001110001110";
            uut_h_1_0 <= "000000000010101110";
            uut_h_0_1 <= "000000000001110101";
            uut_h_1_1 <= "000000010100001001";
            uut_h_0_2 <= "0010111111000101010011";
            uut_h_1_2 <= "0010100101111000101100";
            IF uut_xp_coord /= "0100011100" OR uut_yp_coord /= "0001100011" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1001011";
              state <= "1011101";
            ELSE
              state <= "1010001";
            END IF;
            uut_rst <= '0';
          WHEN "1010001" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0110001110";
            uut_y_coord <= "0110001010";
            uut_h_0_0 <= "000000000100110110";
            uut_h_1_0 <= "000000011011001000";
            uut_h_0_1 <= "000000011001000111";
            uut_h_1_1 <= "000000001000101010";
            uut_h_0_2 <= "0000110110101011001011";
            uut_h_1_2 <= "0001001101000010111010";
            IF uut_xp_coord /= "0110111010" OR uut_yp_coord /= "0111110001" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1001100";
              state <= "1011101";
            ELSE
              state <= "1010010";
            END IF;
            uut_rst <= '0';
          WHEN "1010010" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0101001011";
            uut_y_coord <= "0000111111";
            uut_h_0_0 <= "000000001000111011";
            uut_h_1_0 <= "000000010101100111";
            uut_h_0_1 <= "000000011100111010";
            uut_h_1_1 <= "000000011101000100";
            uut_h_0_2 <= "0010110011010100111100";
            uut_h_1_2 <= "0000111110100001011101";
            IF uut_xp_coord /= "0110111010" OR uut_yp_coord /= "1000011110" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1001101";
              state <= "1011101";
            ELSE
              state <= "1010011";
            END IF;
            uut_rst <= '0';
          WHEN "1010011" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0000010001";
            uut_y_coord <= "0010011100";
            uut_h_0_0 <= "000000001111110000";
            uut_h_1_0 <= "000000010100111101";
            uut_h_0_1 <= "000000011100011110";
            uut_h_1_1 <= "000000010001001110";
            uut_h_0_2 <= "0001000011101110101010";
            uut_h_1_2 <= "0011101010001110101101";
            IF uut_xp_coord /= "1001010001" OR uut_yp_coord /= "0100001100" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1001110";
              state <= "1011101";
            ELSE
              state <= "1010100";
            END IF;
            uut_rst <= '0';
          WHEN "1010100" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0000001111";
            uut_y_coord <= "0110001101";
            uut_h_0_0 <= "000000001111111111";
            uut_h_1_0 <= "000000010011101100";
            uut_h_0_1 <= "000000010010101010";
            uut_h_1_1 <= "000000010110010110";
            uut_h_0_2 <= "0000000111000010100010";
            uut_h_1_2 <= "0001111110101100010001";
            IF uut_xp_coord /= "1011110011" OR uut_yp_coord /= "0110000110" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1001111";
              state <= "1011101";
            ELSE
              state <= "1010101";
            END IF;
            uut_rst <= '0';
          WHEN "1010101" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0010100011";
            uut_y_coord <= "0100000011";
            uut_h_0_0 <= "000101000000000000";
            uut_h_1_0 <= "000000000000000000";
            uut_h_0_1 <= "000000000000000000";
            uut_h_1_1 <= "000101000000000000";
            uut_h_0_2 <= "0000000101011110001100";
            uut_h_1_2 <= "0001100101110001111100";
            IF uut_xp_coord /= "0111100001" OR uut_yp_coord /= "1001110111" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1010000";
              state <= "1011101";
            ELSE
              state <= "1010110";
            END IF;
            uut_rst <= '0';
          WHEN "1010110" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0011001110";
            uut_y_coord <= "0101010001";
            uut_h_0_0 <= "000101000000000000";
            uut_h_1_0 <= "000000000000000000";
            uut_h_0_1 <= "000000000000000000";
            uut_h_1_1 <= "000101000000000000";
            uut_h_0_2 <= "0001110000000001011000";
            uut_h_1_2 <= "0000111100111101100011";
            IF uut_xp_coord /= "0111011110" OR uut_yp_coord /= "1001010110" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1010001";
              state <= "1011101";
            ELSE
              state <= "1010111";
            END IF;
            uut_rst <= '0';
          WHEN "1010111" =>
            uut_input_valid <= '1';
            uut_x_coord <= "0011001010";
            uut_y_coord <= "0000011011";
            uut_h_0_0 <= "000101000000000000";
            uut_h_1_0 <= "000000000000000000";
            uut_h_0_1 <= "000000000000000000";
            uut_h_1_1 <= "000101000000000000";
            uut_h_0_2 <= "0010111001001010000000";
            uut_h_1_2 <= "0010110111100011001000";
            IF uut_xp_coord /= "0111111011" OR uut_yp_coord /= "0110010101" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1010010";
              state <= "1011101";
            ELSE
              state <= "1011000";
            END IF;
            uut_rst <= '0';
          WHEN "1011000" =>
            IF uut_xp_coord /= "0100011010" OR uut_yp_coord /= "1000110011" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1010011";
              state <= "1011101";
            ELSE
              state <= "1011001";
            END IF;
            uut_rst <= '0';
          WHEN "1011001" =>
            IF uut_xp_coord /= "0011111101" OR uut_yp_coord /= "1000011011" OR uut_overflow_x /= '0' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1010100";
              state <= "1011101";
            ELSE
              state <= "1011010";
            END IF;
            uut_rst <= '0';
          WHEN "1011010" =>
            IF uut_overflow_x /= '1' OR uut_overflow_y /= '1' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1010101";
              state <= "1011101";
            ELSE
              state <= "1011011";
            END IF;
            uut_rst <= '0';
          WHEN "1011011" =>
            IF uut_overflow_x /= '1' OR uut_overflow_y /= '1' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1010110";
              state <= "1011101";
            ELSE
              state <= "1011100";
            END IF;
            uut_rst <= '0';
          WHEN "1011100" =>
            IF uut_yp_coord /= "1001111101" OR uut_overflow_x /= '1' OR uut_overflow_y /= '0' OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1010111";
              state <= "1011101";
            ELSE
              state <= "1011101";
            END IF;
            uut_rst <= '0';
          WHEN OTHERS =>
            DONE <= '1';
            uut_rst <= '1';
        END CASE;
      END IF;
    END IF;
  END PROCESS;
END;
