/home/brandyn/fpga-image-registration/modules/./make_a_b_matrices/make_a_b_matrices.vhd