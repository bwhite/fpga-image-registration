/home/brandyn/fpga-image-registration/modules/./convolution/convolution_1x5_gaussian/conv_tb1.vhd