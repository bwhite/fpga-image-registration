/home/brandyn/fpga-image-registration/modules/./pipeline_buffer/pipeline_buffer.vhd