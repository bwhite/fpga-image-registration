/home/brandyn/fpga-image-registration/modules/./image_display_stage/image_display_stage.vhd