/home/brandyn/fpga-image-registration/modules/./smooth_stage/smooth_conv_buffer_3x3.vhd