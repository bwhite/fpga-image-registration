/home/brandyn/fpga-image-registration/modules/./gauss_elim/gauss_elim.vhd