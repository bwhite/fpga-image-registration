/home/brandyn/fpga-image-registration/modules/./smooth_stage/pixel_buffer_3x3.vhd