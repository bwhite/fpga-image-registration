/home/brandyn/fpga-image-registration/modules/./fetch_stage/pixel_conv_buffer.vhd