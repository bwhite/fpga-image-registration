LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
ENTITY make_a_b_matricesT0_tb IS
PORT(
  CLK : IN STD_LOGIC;
  RST : IN STD_LOGIC;
  DONE : OUT STD_LOGIC;
  FAIL : OUT STD_LOGIC;
  FAIL_NUM : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END make_a_b_matricesT0_tb;
ARCHITECTURE behavior OF make_a_b_matricesT0_tb IS
  COMPONENT make_a_b_matrices
  PORT(
    CLK : IN STD_LOGIC;
    RST : IN STD_LOGIC;
    COORD_SHIFT : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    X : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    Y : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    FX : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    FY : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    FT : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    VALID_IN : IN STD_LOGIC;
    DONE : IN STD_LOGIC;
    VALID_OUT : OUT STD_LOGIC;
    DONE_BUF : OUT STD_LOGIC;
    A_0_0 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_0_1 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_0_2 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_0_3 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_0_4 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_0_5 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_1_0 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_1_1 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_1_2 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_1_3 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_1_4 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_1_5 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_2_0 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_2_1 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_2_2 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_2_3 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_2_4 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_2_5 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_3_0 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_3_1 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_3_2 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_3_3 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_3_4 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_3_5 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_4_0 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_4_1 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_4_2 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_4_3 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_4_4 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_4_5 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_5_0 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_5_1 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_5_2 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_5_3 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_5_4 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    A_5_5 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    B_0 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    B_1 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    B_2 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    B_3 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    B_4 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    B_5 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0));
  END COMPONENT;
  SIGNAL uut_rst_wire, uut_rst : STD_LOGIC;
  SIGNAL state : STD_LOGIC_VECTOR(7 DOWNTO 0);
  -- UUT Input
  SIGNAL uut_valid_in, uut_done : STD_LOGIC;
  SIGNAL uut_x, uut_y : STD_LOGIC_VECTOR(11 DOWNTO 0);
  SIGNAL uut_fx, uut_fy, uut_ft : STD_LOGIC_VECTOR(9 DOWNTO 0);
  SIGNAL uut_coord_shift : STD_LOGIC_VECTOR(3 DOWNTO 0);
  -- UUT Output
  SIGNAL uut_valid_out, uut_done_buf : STD_LOGIC;
  SIGNAL uut_a_0_0, uut_a_0_1, uut_a_0_2, uut_a_0_3, uut_a_0_4, uut_a_0_5, uut_a_1_0, uut_a_1_1, uut_a_1_2, uut_a_1_3, uut_a_1_4, uut_a_1_5, uut_a_2_0, uut_a_2_1, uut_a_2_2, uut_a_2_3, uut_a_2_4, uut_a_2_5, uut_a_3_0, uut_a_3_1, uut_a_3_2, uut_a_3_3, uut_a_3_4, uut_a_3_5, uut_a_4_0, uut_a_4_1, uut_a_4_2, uut_a_4_3, uut_a_4_4, uut_a_4_5, uut_a_5_0, uut_a_5_1, uut_a_5_2, uut_a_5_3, uut_a_5_4, uut_a_5_5, uut_b_0, uut_b_1, uut_b_2, uut_b_3, uut_b_4, uut_b_5 : STD_LOGIC_VECTOR(26 DOWNTO 0);
BEGIN
  uut_rst_wire <= RST OR uut_rst;
  uut :  make_a_b_matrices PORT MAP (
    CLK => CLK,
    RST => uut_rst_wire,
    COORD_SHIFT => uut_coord_shift,
    X => uut_x,
    Y => uut_y,
    FX => uut_fx,
    FY => uut_fy,
    FT => uut_ft,
    VALID_IN => uut_valid_in,
    DONE => uut_done,
    VALID_OUT => uut_valid_out,
    DONE_BUF => uut_done_buf,
    A_0_0 => uut_a_0_0,
    A_0_1 => uut_a_0_1,
    A_0_2 => uut_a_0_2,
    A_0_3 => uut_a_0_3,
    A_0_4 => uut_a_0_4,
    A_0_5 => uut_a_0_5,
    A_1_0 => uut_a_1_0,
    A_1_1 => uut_a_1_1,
    A_1_2 => uut_a_1_2,
    A_1_3 => uut_a_1_3,
    A_1_4 => uut_a_1_4,
    A_1_5 => uut_a_1_5,
    A_2_0 => uut_a_2_0,
    A_2_1 => uut_a_2_1,
    A_2_2 => uut_a_2_2,
    A_2_3 => uut_a_2_3,
    A_2_4 => uut_a_2_4,
    A_2_5 => uut_a_2_5,
    A_3_0 => uut_a_3_0,
    A_3_1 => uut_a_3_1,
    A_3_2 => uut_a_3_2,
    A_3_3 => uut_a_3_3,
    A_3_4 => uut_a_3_4,
    A_3_5 => uut_a_3_5,
    A_4_0 => uut_a_4_0,
    A_4_1 => uut_a_4_1,
    A_4_2 => uut_a_4_2,
    A_4_3 => uut_a_4_3,
    A_4_4 => uut_a_4_4,
    A_4_5 => uut_a_4_5,
    A_5_0 => uut_a_5_0,
    A_5_1 => uut_a_5_1,
    A_5_2 => uut_a_5_2,
    A_5_3 => uut_a_5_3,
    A_5_4 => uut_a_5_4,
    A_5_5 => uut_a_5_5,
    B_0 => uut_b_0,
    B_1 => uut_b_1,
    B_2 => uut_b_2,
    B_3 => uut_b_3,
    B_4 => uut_b_4,
    B_5 => uut_b_5
  );
  PROCESS (CLK) IS
  BEGIN
    IF CLK'event AND CLK='1' THEN
      IF RST='1' THEN
        DONE <= '0';
        FAIL <= '0';
        uut_rst <= '1';
        FAIL_NUM <= (OTHERS => '0');
        state <= (OTHERS => '0');
      ELSE
        CASE state IS
          WHEN "00000000" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000101100";
            uut_y <= "000000000111";
            uut_fx <= "0110111000";
            uut_fy <= "0011001001";
            uut_ft <= "0001010101";
            uut_valid_in <= '1';
            uut_done <= '0';
            state <= "00000001";
            uut_rst <= '0';
          WHEN "00000001" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000101000";
            uut_y <= "000000110000";
            uut_fx <= "0111110101";
            uut_fy <= "1000000001";
            uut_ft <= "0101110110";
            uut_valid_in <= '1';
            uut_done <= '0';
            state <= "00000010";
            uut_rst <= '0';
          WHEN "00000010" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000001110";
            uut_y <= "000000111110";
            uut_fx <= "0000011100";
            uut_fy <= "1111101011";
            uut_ft <= "0100110101";
            uut_valid_in <= '1';
            uut_done <= '0';
            state <= "00000011";
            uut_rst <= '0';
          WHEN "00000011" =>
            uut_coord_shift <= "0101";
            uut_x <= "111111011110";
            uut_y <= "000000000000";
            uut_fx <= "0110011010";
            uut_fy <= "0001001100";
            uut_ft <= "0101100001";
            uut_valid_in <= '1';
            uut_done <= '0';
            state <= "00000100";
            uut_rst <= '0';
          WHEN "00000100" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000011110";
            uut_y <= "000000001011";
            uut_fx <= "1011111101";
            uut_fy <= "0010101010";
            uut_ft <= "1001010101";
            uut_valid_in <= '1';
            uut_done <= '0';
            state <= "00000101";
            uut_rst <= '0';
          WHEN "00000101" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000010000";
            uut_y <= "000000010100";
            uut_fx <= "0011101011";
            uut_fy <= "0110010000";
            uut_ft <= "0111101110";
            uut_valid_in <= '1';
            uut_done <= '0';
            state <= "00000110";
            uut_rst <= '0';
          WHEN "00000110" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000100010";
            uut_y <= "000000001010";
            uut_fx <= "0110110111";
            uut_fy <= "0001010010";
            uut_ft <= "1000010001";
            uut_valid_in <= '1';
            uut_done <= '0';
            state <= "00000111";
            uut_rst <= '0';
          WHEN "00000111" =>
            uut_coord_shift <= "0101";
            uut_x <= "111111010000";
            uut_y <= "000000101110";
            uut_fx <= "1111110000";
            uut_fy <= "0101100001";
            uut_ft <= "1011010110";
            uut_valid_in <= '1';
            uut_done <= '0';
            state <= "00001000";
            uut_rst <= '0';
          WHEN "00001000" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000000110";
            uut_y <= "000000010000";
            uut_fx <= "1000100001";
            uut_fy <= "0001110101";
            uut_ft <= "1101110011";
            uut_valid_in <= '1';
            uut_done <= '0';
            state <= "00001001";
            uut_rst <= '0';
          WHEN "00001001" =>
            uut_coord_shift <= "0101";
            uut_x <= "111111000111";
            uut_y <= "111111111111";
            uut_fx <= "1011000101";
            uut_fy <= "1001111110";
            uut_ft <= "1011010010";
            uut_valid_in <= '1';
            uut_done <= '0';
            state <= "00001010";
            uut_rst <= '0';
          WHEN "00001010" =>
            uut_coord_shift <= "0101";
            uut_x <= "111111010011";
            uut_y <= "111111011001";
            uut_fx <= "1000101100";
            uut_fy <= "0010001010";
            uut_ft <= "1100100001";
            uut_valid_in <= '1';
            uut_done <= '0';
            state <= "00001011";
            uut_rst <= '0';
          WHEN "00001011" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000000100";
            uut_y <= "000000011000";
            uut_fx <= "1111111111";
            uut_fy <= "0000100101";
            uut_ft <= "1111001000";
            uut_valid_in <= '1';
            uut_done <= '0';
            state <= "00001100";
            uut_rst <= '0';
          WHEN "00001100" =>
            uut_coord_shift <= "0101";
            uut_x <= "111111010000";
            uut_y <= "111111111111";
            uut_fx <= "0101101001";
            uut_fy <= "0101111111";
            uut_ft <= "1100010101";
            uut_valid_in <= '1';
            uut_done <= '0';
            state <= "00001101";
            uut_rst <= '0';
          WHEN "00001101" =>
            uut_coord_shift <= "0101";
            uut_x <= "111111011011";
            uut_y <= "000000001000";
            uut_fx <= "0010010000";
            uut_fy <= "1110101011";
            uut_ft <= "1011010011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000101111010001000000000" OR uut_a_0_1 /= "010000001111110110000000000" OR uut_a_0_2 /= "000010100101011011100000000" OR uut_a_0_3 /= "000000010101100101111000000" OR uut_a_0_4 /= "000111011011000001010000000" OR uut_a_0_5 /= "000001001011100100100100000" OR uut_a_1_0 /= "000000100000011111101100000" OR uut_a_1_1 /= "001011001010111001001000000" OR uut_a_1_2 /= "000001110001101110111010000" OR uut_a_1_3 /= "000000001110110110000010100" OR uut_a_1_4 /= "000101000110100100110111000" OR uut_a_1_5 /= "000000110011111101001000110" OR uut_a_2_0 /= "000000000101001010110111000" OR uut_a_2_1 /= "000001110001101110111010000" OR uut_a_2_2 /= "000000010010000110000000100" OR uut_a_2_3 /= "000000000010010111001001001" OR uut_a_2_4 /= "000000110011111101001000110" OR uut_a_2_5 /= "000000001000010000111111111" OR uut_a_3_0 /= "000000010101100101111000000" OR uut_a_3_1 /= "000111011011000001010000000" OR uut_a_3_2 /= "000001001011100100100100000" OR uut_a_3_3 /= "000000001001110111010001000" OR uut_a_3_4 /= "000011011000111111110110000" OR uut_a_3_5 /= "000000100010100001011011100" OR uut_a_4_0 /= "000000001110110110000010100" OR uut_a_4_1 /= "000101000110100100110111000" OR uut_a_4_2 /= "000000110011111101001000110" OR uut_a_4_3 /= "000000000110110001111111101" OR uut_a_4_4 /= "000010010101001011111001001" OR uut_a_4_5 /= "000000010111101110111110111" OR uut_a_5_0 /= "000000000010010111001001001" OR uut_a_5_1 /= "000000110011111101001000110" OR uut_a_5_2 /= "000000001000010000111111111" OR uut_a_5_3 /= "000000000001000101000010110" OR uut_a_5_4 /= "000000010111101110111110111" OR uut_a_5_5 /= "000000000011110001101010000" THEN
              FAIL <= '1';
              FAIL_NUM <= "00000000";
              state <= "11111101";
            ELSE
              state <= "00001110";
            END IF;
            uut_rst <= '0';
          WHEN "00001110" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000111001";
            uut_y <= "111111001011";
            uut_fx <= "1001101100";
            uut_fy <= "1010010001";
            uut_ft <= "1010101010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000111101010001111001000" OR uut_a_0_1 /= "010011001001100101110100000" OR uut_a_0_2 /= "010110111110101101011000000" OR uut_a_0_3 /= "111111000001011111110101000" OR uut_a_0_4 /= "101100011101111100100100000" OR uut_a_0_5 /= "101000100011111011111000000" OR uut_a_1_0 /= "000000100110010011001011101" OR uut_a_1_1 /= "001011111101111111101000100" OR uut_a_1_2 /= "001110010111001100010111000" OR uut_a_1_3 /= "111111011000111011111001001" OR uut_a_1_4 /= "110011110010101101110110100" OR uut_a_1_5 /= "110001010110011101011011000" OR uut_a_2_0 /= "000000101101111101011010110" OR uut_a_2_1 /= "001110010111001100010111000" OR uut_a_2_2 /= "010001001111000010000010000" OR uut_a_2_3 /= "111111010001000111110111110" OR uut_a_2_4 /= "110001010110011101011011000" OR uut_a_2_5 /= "101110011010111100111010000" OR uut_a_3_0 /= "111111000001011111110101000" OR uut_a_3_1 /= "101100011101111100100100000" OR uut_a_3_2 /= "101000100011111011111000000" OR uut_a_3_3 /= "000000111111110000000001000" OR uut_a_3_4 /= "010011111011000000010100000" OR uut_a_3_5 /= "010111111010000000011000000" OR uut_a_4_0 /= "111111011000111011111001001" OR uut_a_4_1 /= "110011110010101101110110100" OR uut_a_4_2 /= "110001010110011101011011000" OR uut_a_4_3 /= "000000100111110110000000101" OR uut_a_4_4 /= "001100011100111000001100100" OR uut_a_4_5 /= "001110111100010000001111000" OR uut_a_5_0 /= "111111010001000111110111110" OR uut_a_5_1 /= "110001010110011101011011000" OR uut_a_5_2 /= "101110011010111100111010000" OR uut_a_5_3 /= "000000101111110100000000110" OR uut_a_5_4 /= "001110111100010000001111000" OR uut_a_5_5 /= "010001111011100000010010000" THEN
              FAIL <= '1';
              FAIL_NUM <= "00000001";
              state <= "11111101";
            ELSE
              state <= "00001111";
            END IF;
            uut_rst <= '0';
          WHEN "00001111" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000001111";
            uut_y <= "000000001001";
            uut_fx <= "1000110101";
            uut_fy <= "0110111010";
            uut_ft <= "0011101010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000001100010000000" OR uut_a_0_1 /= "000000000001010101110000000" OR uut_a_0_2 /= "000000000101111011110000000" OR uut_a_0_3 /= "111111111111110110110100000" OR uut_a_0_4 /= "111111111110111111101100000" OR uut_a_0_5 /= "111111111011100011001100000" OR uut_a_1_0 /= "000000000000000010101011100" OR uut_a_1_1 /= "000000000000010010110000100" OR uut_a_1_2 /= "000000000001010011000100100" OR uut_a_1_3 /= "111111111111111101111111011" OR uut_a_1_4 /= "111111111111110001111011101" OR uut_a_1_5 /= "111111111111000001101100101" OR uut_a_2_0 /= "000000000000001011110111100" OR uut_a_2_1 /= "000000000001010011000100100" OR uut_a_2_2 /= "000000000101101111111000100" OR uut_a_2_3 /= "111111111111110111000110011" OR uut_a_2_4 /= "111111111111000001101100101" OR uut_a_2_5 /= "111111111011101100000101101" OR uut_a_3_0 /= "111111111111110110110100000" OR uut_a_3_1 /= "111111111110111111101100000" OR uut_a_3_2 /= "111111111011100011001100000" OR uut_a_3_3 /= "000000000000000110111001000" OR uut_a_3_4 /= "000000000000110000001111000" OR uut_a_3_5 /= "000000000011010101100111000" OR uut_a_4_0 /= "111111111111111101111111011" OR uut_a_4_1 /= "111111111111110001111011101" OR uut_a_4_2 /= "111111111111000001101100101" OR uut_a_4_3 /= "000000000000000001100000011" OR uut_a_4_4 /= "000000000000001010100011010" OR uut_a_4_5 /= "000000000000101110101110100" OR uut_a_5_0 /= "111111111111110111000110011" OR uut_a_5_1 /= "111111111111000001101100101" OR uut_a_5_2 /= "111111111011101100000101101" OR uut_a_5_3 /= "000000000000000110101011001" OR uut_a_5_4 /= "000000000000101110101110100" OR uut_a_5_5 /= "000000000011001110111011110" THEN
              FAIL <= '1';
              FAIL_NUM <= "00000010";
              state <= "11111101";
            ELSE
              state <= "00010000";
            END IF;
            uut_rst <= '0';
          WHEN "00010000" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000011110";
            uut_y <= "111111001001";
            uut_fx <= "0101110001";
            uut_fy <= "0110111101";
            uut_ft <= "0111110000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000101001000010100100000" OR uut_a_0_1 /= "110101000110010100011100000" OR uut_a_0_2 /= "000000000000000000000000000" OR uut_a_0_3 /= "000000000111100110111000000" OR uut_a_0_4 /= "111101111110101011001000000" OR uut_a_0_5 /= "000000000000000000000000000" OR uut_a_1_0 /= "111111101010001100101000111" OR uut_a_1_1 /= "000101110010101001001001001" OR uut_a_1_2 /= "000000000000000000000000000" OR uut_a_1_3 /= "111111111011111101010110010" OR uut_a_1_4 /= "000001000100101101000101110" OR uut_a_1_5 /= "000000000000000000000000000" OR uut_a_2_0 /= "000000000000000000000000000" OR uut_a_2_1 /= "000000000000000000000000000" OR uut_a_2_2 /= "000000000000000000000000000" OR uut_a_2_3 /= "000000000000000000000000000" OR uut_a_2_4 /= "000000000000000000000000000" OR uut_a_2_5 /= "000000000000000000000000000" OR uut_a_3_0 /= "000000000111100110111000000" OR uut_a_3_1 /= "111101111110101011001000000" OR uut_a_3_2 /= "000000000000000000000000000" OR uut_a_3_3 /= "000000000001011010010000000" OR uut_a_3_4 /= "111111101000000001110000000" OR uut_a_3_5 /= "000000000000000000000000000" OR uut_a_4_0 /= "111111111011111101010110010" OR uut_a_4_1 /= "000001000100101101000101110" OR uut_a_4_2 /= "000000000000000000000000000" OR uut_a_4_3 /= "111111111111010000000011100" OR uut_a_4_4 /= "000000001100101111000100100" OR uut_a_4_5 /= "000000000000000000000000000" OR uut_a_5_0 /= "000000000000000000000000000" OR uut_a_5_1 /= "000000000000000000000000000" OR uut_a_5_2 /= "000000000000000000000000000" OR uut_a_5_3 /= "000000000000000000000000000" OR uut_a_5_4 /= "000000000000000000000000000" OR uut_a_5_5 /= "000000000000000000000000000" THEN
              FAIL <= '1';
              FAIL_NUM <= "00000011";
              state <= "11111101";
            ELSE
              state <= "00010001";
            END IF;
            uut_rst <= '0';
          WHEN "00010001" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000101101";
            uut_y <= "000000100100";
            uut_fx <= "0000001110";
            uut_fy <= "1010110110";
            uut_ft <= "1110011000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000010000011000001001000" OR uut_a_0_1 /= "000011110101101010000111000" OR uut_a_0_2 /= "000001011010000100110001100" OR uut_a_0_3 /= "111111110101010000000010000" OR uut_a_0_4 /= "111101011110110000011110000" OR uut_a_0_5 /= "111111000100111000001011000" OR uut_a_1_0 /= "000000000111101011010100001" OR uut_a_1_1 /= "000001110011001001101111010" OR uut_a_1_2 /= "000000101010001110001111001" OR uut_a_1_3 /= "111111111010111101100000111" OR uut_a_1_4 /= "111110110100011010101110000" OR uut_a_1_5 /= "111111100100010010010101001" OR uut_a_2_0 /= "000000000010110100001001100" OR uut_a_2_1 /= "000000101010001110001111001" OR uut_a_2_2 /= "000000001111011110110100100" OR uut_a_2_3 /= "111111111110001001110000010" OR uut_a_2_4 /= "111111100100010010010101001" OR uut_a_2_5 /= "111111110101110101101001111" OR uut_a_3_0 /= "111111110101010000000010000" OR uut_a_3_1 /= "111101011110110000011110000" OR uut_a_3_2 /= "111111000100111000001011000" OR uut_a_3_3 /= "000000000111000011100100000" OR uut_a_3_4 /= "000001101001110101011100000" OR uut_a_3_5 /= "000000100110110011100110000" OR uut_a_4_0 /= "111111111010111101100000111" OR uut_a_4_1 /= "111110110100011010101110000" OR uut_a_4_2 /= "111111100100010010010101001" OR uut_a_4_3 /= "000000000011010011101010111" OR uut_a_4_4 /= "000000110001100111000011001" OR uut_a_4_5 /= "000000010010001100001011110" OR uut_a_5_0 /= "111111111110001001110000010" OR uut_a_5_1 /= "111111100100010010010101001" OR uut_a_5_2 /= "111111110101110101101001111" OR uut_a_5_3 /= "000000000001001101100111001" OR uut_a_5_4 /= "000000010010001100001011110" OR uut_a_5_5 /= "000000000110101010110111100" THEN
              FAIL <= '1';
              FAIL_NUM <= "00000100";
              state <= "11111101";
            ELSE
              state <= "00010010";
            END IF;
            uut_rst <= '0';
          WHEN "00010010" =>
            uut_coord_shift <= "0101";
            uut_x <= "111111010010";
            uut_y <= "111111000100";
            uut_fx <= "0111000010";
            uut_fy <= "1100110101";
            uut_ft <= "1100101111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000001101011110111001000" OR uut_a_0_1 /= "000001101011110111001000000" OR uut_a_0_2 /= "000010000110110100111010000" OR uut_a_0_3 /= "000000010110111100110000000" OR uut_a_0_4 /= "000010110111100110000000000" OR uut_a_0_5 /= "000011100101011111100000000" OR uut_a_1_0 /= "000000000011010111101110010" OR uut_a_1_1 /= "000000011010111101110010000" OR uut_a_1_2 /= "000000100001101101001110100" OR uut_a_1_3 /= "000000000101101111001100000" OR uut_a_1_4 /= "000000101101111001100000000" OR uut_a_1_5 /= "000000111001010111111000000" OR uut_a_2_0 /= "000000000100001101101001110" OR uut_a_2_1 /= "000000100001101101001110100" OR uut_a_2_2 /= "000000101010001000100010001" OR uut_a_2_3 /= "000000000111001010111111000" OR uut_a_2_4 /= "000000111001010111111000000" OR uut_a_2_5 /= "000001000111101101110110000" OR uut_a_3_0 /= "000000010110111100110000000" OR uut_a_3_1 /= "000010110111100110000000000" OR uut_a_3_2 /= "000011100101011111100000000" OR uut_a_3_3 /= "000000100111000100000000000" OR uut_a_3_4 /= "000100111000100000000000000" OR uut_a_3_5 /= "000110000110101000000000000" OR uut_a_4_0 /= "000000000101101111001100000" OR uut_a_4_1 /= "000000101101111001100000000" OR uut_a_4_2 /= "000000111001010111111000000" OR uut_a_4_3 /= "000000001001110001000000000" OR uut_a_4_4 /= "000001001110001000000000000" OR uut_a_4_5 /= "000001100001101010000000000" OR uut_a_5_0 /= "000000000111001010111111000" OR uut_a_5_1 /= "000000111001010111111000000" OR uut_a_5_2 /= "000001000111101101110110000" OR uut_a_5_3 /= "000000001100001101010000000" OR uut_a_5_4 /= "000001100001101010000000000" OR uut_a_5_5 /= "000001111010000100100000000" THEN
              FAIL <= '1';
              FAIL_NUM <= "00000101";
              state <= "11111101";
            ELSE
              state <= "00010011";
            END IF;
            uut_rst <= '0';
          WHEN "00010011" =>
            uut_coord_shift <= "0101";
            uut_x <= "111111101011";
            uut_y <= "111111111100";
            uut_fx <= "0010011000";
            uut_fy <= "1000011010";
            uut_ft <= "0101011110";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000101111000011010001000" OR uut_a_0_1 /= "001100011111110111100001000" OR uut_a_0_2 /= "000011101011010000010101000" OR uut_a_0_3 /= "000000001000110010011110000" OR uut_a_0_4 /= "000010010101011001111110000" OR uut_a_0_5 /= "000000101011111100010110000" OR uut_a_1_0 /= "000000011000111111101111000" OR uut_a_1_1 /= "000110101000111011011111100" OR uut_a_1_2 /= "000001111100111110101011001" OR uut_a_1_3 /= "000000000100101010110011111" OR uut_a_1_4 /= "000001001111010111110010111" OR uut_a_1_5 /= "000000010111010110000011101" OR uut_a_2_0 /= "000000000111010110100000101" OR uut_a_2_1 /= "000001111100111110101011001" OR uut_a_2_2 /= "000000100100110000100011010" OR uut_a_2_3 /= "000000000001010111111000101" OR uut_a_2_4 /= "000000010111010110000011101" OR uut_a_2_5 /= "000000000110110111011011011" OR uut_a_3_0 /= "000000001000110010011110000" OR uut_a_3_1 /= "000010010101011001111110000" OR uut_a_3_2 /= "000000101011111100010110000" OR uut_a_3_3 /= "000000000001101001000100000" OR uut_a_3_4 /= "000000011011111010000100000" OR uut_a_3_5 /= "000000001000001101010100000" OR uut_a_4_0 /= "000000000100101010110011111" OR uut_a_4_1 /= "000001001111010111110010111" OR uut_a_4_2 /= "000000010111010110000011101" OR uut_a_4_3 /= "000000000000110111110100001" OR uut_a_4_4 /= "000000001110110100110110001" OR uut_a_4_5 /= "000000000100010111000100101" OR uut_a_5_0 /= "000000000001010111111000101" OR uut_a_5_1 /= "000000010111010110000011101" OR uut_a_5_2 /= "000000000110110111011011011" OR uut_a_5_3 /= "000000000000010000011010101" OR uut_a_5_4 /= "000000000100010111000100101" OR uut_a_5_5 /= "000000000001010010000101001" THEN
              FAIL <= '1';
              FAIL_NUM <= "00000110";
              state <= "11111101";
            ELSE
              state <= "00010100";
            END IF;
            uut_rst <= '0';
          WHEN "00010100" =>
            uut_coord_shift <= "0110";
            uut_x <= "000000001111";
            uut_y <= "000001011010";
            uut_fx <= "1101100100";
            uut_fy <= "1111001001";
            uut_ft <= "1000111000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000100000000000" OR uut_a_0_1 /= "111111111110100000000000000" OR uut_a_0_2 /= "000000000001011100000000000" OR uut_a_0_3 /= "111111111110100111110000000" OR uut_a_0_4 /= "000000100001000110000000000" OR uut_a_0_5 /= "111111100000010010010000000" OR uut_a_1_0 /= "111111111111111101000000000" OR uut_a_1_1 /= "000000000001001000000000000" OR uut_a_1_2 /= "111111111110111011000000000" OR uut_a_1_3 /= "000000000001000010001100000" OR uut_a_1_4 /= "111111100111001011100000000" OR uut_a_1_5 /= "000000010111110010010100000" OR uut_a_2_0 /= "000000000000000010111000000" OR uut_a_2_1 /= "111111111110111011000000000" OR uut_a_2_2 /= "000000000001000010001000000" OR uut_a_2_3 /= "111111111111000000100100100" OR uut_a_2_4 /= "000000010111110010010100000" OR uut_a_2_5 /= "111111101001001101000111100" OR uut_a_3_0 /= "111111111110100111110000000" OR uut_a_3_1 /= "000000100001000110000000000" OR uut_a_3_2 /= "111111100000010010010000000" OR uut_a_3_3 /= "000000011110011011000001000" OR uut_a_3_4 /= "110100100101110111101000000" OR uut_a_3_5 /= "001010111011101101010111000" OR uut_a_4_0 /= "000000000001000010001100000" OR uut_a_4_1 /= "111111100111001011100000000" OR uut_a_4_2 /= "000000010111110010010100000" OR uut_a_4_3 /= "111111101001001011101111010" OR uut_a_4_4 /= "001000100011100110010010000" OR uut_a_4_5 /= "110111110011001101111110110" OR uut_a_5_0 /= "111111111111000000100100100" OR uut_a_5_1 /= "000000010111110010010100000" OR uut_a_5_2 /= "111111101001001101000111100" OR uut_a_5_3 /= "000000010101110111011010101" OR uut_a_5_4 /= "110111110011001101111110110" OR uut_a_5_5 /= "000111110110111010100110100" THEN
              FAIL <= '1';
              FAIL_NUM <= "00000111";
              state <= "11111101";
            ELSE
              state <= "00010101";
            END IF;
            uut_rst <= '0';
          WHEN "00010101" =>
            uut_coord_shift <= "0110";
            uut_x <= "111110101110";
            uut_y <= "000000101001";
            uut_fx <= "1101010011";
            uut_fy <= "0110011000";
            uut_ft <= "1001111001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000111000000001000001000" OR uut_a_0_1 /= "000010101000000011000011000" OR uut_a_0_2 /= "000111000000001000001000000" OR uut_a_0_3 /= "111111110010010100010101000" OR uut_a_0_4 /= "111111010110111100111111000" OR uut_a_0_5 /= "111110010010100010101000000" OR uut_a_1_0 /= "000000000101010000000110000" OR uut_a_1_1 /= "000000001111110000010010010" OR uut_a_1_2 /= "000000101010000000110000110" OR uut_a_1_3 /= "111111111110101101111001111" OR uut_a_1_4 /= "111111111100001001101101111" OR uut_a_1_5 /= "111111110101101111001111110" OR uut_a_2_0 /= "000000001110000000010000010" OR uut_a_2_1 /= "000000101010000000110000110" OR uut_a_2_2 /= "000001110000000010000010000" OR uut_a_2_3 /= "111111111100100101000101010" OR uut_a_2_4 /= "111111110101101111001111110" OR uut_a_2_5 /= "111111100100101000101010000" OR uut_a_3_0 /= "111111110010010100010101000" OR uut_a_3_1 /= "111111010110111100111111000" OR uut_a_3_2 /= "111110010010100010101000000" OR uut_a_3_3 /= "000000000011010101111001000" OR uut_a_3_4 /= "000000001010000001101011000" OR uut_a_3_5 /= "000000011010101111001000000" OR uut_a_4_0 /= "111111111110101101111001111" OR uut_a_4_1 /= "111111111100001001101101111" OR uut_a_4_2 /= "111111110101101111001111110" OR uut_a_4_3 /= "000000000000010100000011010" OR uut_a_4_4 /= "000000000000111100001010000" OR uut_a_4_5 /= "000000000010100000011010110" OR uut_a_5_0 /= "111111111100100101000101010" OR uut_a_5_1 /= "111111110101101111001111110" OR uut_a_5_2 /= "111111100100101000101010000" OR uut_a_5_3 /= "000000000000110101011110010" OR uut_a_5_4 /= "000000000010100000011010110" OR uut_a_5_5 /= "000000000110101011110010000" THEN
              FAIL <= '1';
              FAIL_NUM <= "00001000";
              state <= "11111101";
            ELSE
              state <= "00010110";
            END IF;
            uut_rst <= '0';
          WHEN "00010110" =>
            uut_coord_shift <= "0110";
            uut_x <= "000001111101";
            uut_y <= "000000001010";
            uut_fx <= "0011010100";
            uut_fy <= "0111111111";
            uut_ft <= "1100100111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000011000001110011001000" OR uut_a_0_1 /= "110101001101100101110111100" OR uut_a_0_2 /= "111111110011111000110011100" OR uut_a_0_3 /= "000000011101101011110110000" OR uut_a_0_4 /= "110010110001111110011101000" OR uut_a_0_5 /= "111111110001001010000101000" OR uut_a_1_0 /= "111111101010011011001011101" OR uut_a_1_1 /= "001001100110111001010001100" OR uut_a_1_2 /= "000000001010110010011010001" OR uut_a_1_3 /= "111111100101100011111100111" OR uut_a_1_4 /= "001011110001011111011000001" OR uut_a_1_5 /= "000000001101001110000001100" OR uut_a_2_0 /= "111111111111100111110001100" OR uut_a_2_1 /= "000000001010110010011010001" OR uut_a_2_2 /= "000000000000001100000111001" OR uut_a_2_3 /= "111111111111100010010100001" OR uut_a_2_4 /= "000000001101001110000001100" OR uut_a_2_5 /= "000000000000001110110101111" OR uut_a_3_0 /= "000000011101101011110110000" OR uut_a_3_1 /= "110010110001111110011101000" OR uut_a_3_2 /= "111111110001001010000101000" OR uut_a_3_3 /= "000000100100011000000100000" OR uut_a_3_4 /= "101111110011010010001110000" OR uut_a_3_5 /= "111111101101110011111110000" OR uut_a_4_0 /= "111111100101100011111100111" OR uut_a_4_1 /= "001011110001011111011000001" OR uut_a_4_2 /= "000000001101001110000001100" OR uut_a_4_3 /= "111111011111100110100100011" OR uut_a_4_4 /= "001110011011010100110001100" OR uut_a_4_5 /= "000000010000001100101101110" OR uut_a_5_0 /= "111111111111100010010100001" OR uut_a_5_1 /= "000000001101001110000001100" OR uut_a_5_2 /= "000000000000001110110101111" OR uut_a_5_3 /= "111111111111011011100111111" OR uut_a_5_4 /= "000000010000001100101101110" OR uut_a_5_5 /= "000000000000010010001100000" THEN
              FAIL <= '1';
              FAIL_NUM <= "00001001";
              state <= "11111101";
            ELSE
              state <= "00010111";
            END IF;
            uut_rst <= '0';
          WHEN "00010111" =>
            uut_coord_shift <= "0110";
            uut_x <= "111111101011";
            uut_y <= "111111110111";
            uut_fx <= "0100001110";
            uut_fy <= "0101000110";
            uut_ft <= "1001100111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000110101011110010000000" OR uut_a_0_1 /= "101101001100110111011000000" OR uut_a_0_2 /= "101111101101010010001000000" OR uut_a_0_3 /= "111111110000001110111000000" OR uut_a_0_4 /= "000101100010110001010100000" OR uut_a_0_5 /= "000100110011011101111100000" OR uut_a_1_0 /= "111111011010011001101110110" OR uut_a_1_1 /= "001101001101111101000100001" OR uut_a_1_2 /= "001011011101001010010000011" OR uut_a_1_3 /= "000000001011000101100010101" OR uut_a_1_4 /= "111100000110100011010100111" OR uut_a_1_5 /= "111100100111110011111100110" OR uut_a_2_0 /= "111111011111011010100100010" OR uut_a_2_1 /= "001011011101001010010000011" OR uut_a_2_2 /= "001001111011011001111101001" OR uut_a_2_3 /= "000000001001100110111011111" OR uut_a_2_4 /= "111100100111110011111100110" OR uut_a_2_5 /= "111101000100101000110000011" OR uut_a_3_0 /= "111111110000001110111000000" OR uut_a_3_1 /= "000101100010110001010100000" OR uut_a_3_2 /= "000100110011011101111100000" OR uut_a_3_3 /= "000000000100101001100100000" OR uut_a_3_4 /= "111110010111011000110110000" OR uut_a_3_5 /= "111110100101010101100010000" OR uut_a_4_0 /= "000000001011000101100010101" OR uut_a_4_1 /= "111100000110100011010100111" OR uut_a_4_2 /= "111100100111110011111100110" OR uut_a_4_3 /= "111111111100101110110001101" OR uut_a_4_4 /= "000001001001100011100010000" OR uut_a_4_5 /= "000000111111101111110111000" OR uut_a_5_0 /= "000000001001100110111011111" OR uut_a_5_1 /= "111100100111110011111100110" OR uut_a_5_2 /= "111101000100101000110000011" OR uut_a_5_3 /= "111111111101001010101011000" OR uut_a_5_4 /= "000000111111101111110111000" OR uut_a_5_5 /= "000000110111001111111000010" THEN
              FAIL <= '1';
              FAIL_NUM <= "00001010";
              state <= "11111101";
            ELSE
              state <= "00011000";
            END IF;
            uut_rst <= '0';
          WHEN "00011000" =>
            uut_coord_shift <= "0110";
            uut_x <= "111110101110";
            uut_y <= "111111011101";
            uut_fx <= "1000111010";
            uut_fy <= "0000010110";
            uut_ft <= "1101011000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000000000001000" OR uut_a_0_1 /= "000000000000000000000010000" OR uut_a_0_2 /= "000000000000000000001100000" OR uut_a_0_3 /= "111111111111111111011011000" OR uut_a_0_4 /= "111111111111111110110110000" OR uut_a_0_5 /= "111111111111111001000100000" OR uut_a_1_0 /= "000000000000000000000000000" OR uut_a_1_1 /= "000000000000000000000000001" OR uut_a_1_2 /= "000000000000000000000000110" OR uut_a_1_3 /= "111111111111111111111101101" OR uut_a_1_4 /= "111111111111111111111011011" OR uut_a_1_5 /= "111111111111111111100100010" OR uut_a_2_0 /= "000000000000000000000000011" OR uut_a_2_1 /= "000000000000000000000000110" OR uut_a_2_2 /= "000000000000000000000100100" OR uut_a_2_3 /= "111111111111111111110010001" OR uut_a_2_4 /= "111111111111111111100100010" OR uut_a_2_5 /= "111111111111111101011001100" OR uut_a_3_0 /= "111111111111111111011011000" OR uut_a_3_1 /= "111111111111111110110110000" OR uut_a_3_2 /= "111111111111111001000100000" OR uut_a_3_3 /= "000000000000010101011001000" OR uut_a_3_4 /= "000000000000101010110010000" OR uut_a_3_5 /= "000000000100000000101100000" OR uut_a_4_0 /= "111111111111111111111101101" OR uut_a_4_1 /= "111111111111111111111011011" OR uut_a_4_2 /= "111111111111111111100100010" OR uut_a_4_3 /= "000000000000000001010101100" OR uut_a_4_4 /= "000000000000000010101011001" OR uut_a_4_5 /= "000000000000010000000010110" OR uut_a_5_0 /= "111111111111111111110010001" OR uut_a_5_1 /= "111111111111111111100100010" OR uut_a_5_2 /= "111111111111111101011001100" OR uut_a_5_3 /= "000000000000001000000001011" OR uut_a_5_4 /= "000000000000010000000010110" OR uut_a_5_5 /= "000000000001100000010000100" THEN
              FAIL <= '1';
              FAIL_NUM <= "00001011";
              state <= "11111101";
            ELSE
              state <= "00011001";
            END IF;
            uut_rst <= '0';
          WHEN "00011001" =>
            uut_coord_shift <= "0110";
            uut_x <= "111110101101";
            uut_y <= "111110110110";
            uut_fx <= "0110011111";
            uut_fy <= "0010110100";
            uut_ft <= "1111100000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000011111110100010001000" OR uut_a_0_1 /= "110100000100011001101000000" OR uut_a_0_2 /= "111111110000000101110111100" OR uut_a_0_3 /= "000000100001110000010111000" OR uut_a_0_4 /= "110011010101110111011000000" OR uut_a_0_5 /= "111111101111000111110100100" OR uut_a_1_0 /= "111111101000001000110011010" OR uut_a_1_1 /= "001000111100101100110010000" OR uut_a_1_2 /= "000000001011111011100110011" OR uut_a_1_3 /= "111111100110101011101110110" OR uut_a_1_4 /= "001001011111100110011110000" OR uut_a_1_5 /= "000000001100101010001000101" OR uut_a_2_0 /= "111111111111100000001011101" OR uut_a_2_1 /= "000000001011111011100110011" OR uut_a_2_2 /= "000000000000001111111010001" OR uut_a_2_3 /= "111111111111011110001111101" OR uut_a_2_4 /= "000000001100101010001000101" OR uut_a_2_5 /= "000000000000010000111000001" OR uut_a_3_0 /= "000000100001110000010111000" OR uut_a_3_1 /= "110011010101110111011000000" OR uut_a_3_2 /= "111111101111000111110100100" OR uut_a_3_3 /= "000000100011110100000001000" OR uut_a_3_4 /= "110010100100011111101000000" OR uut_a_3_5 /= "111111101110000101111111100" OR uut_a_4_0 /= "111111100110101011101110110" OR uut_a_4_1 /= "001001011111100110011110000" OR uut_a_4_2 /= "000000001100101010001000101" OR uut_a_4_3 /= "111111100101001000111111010" OR uut_a_4_4 /= "001010000100101000010010000" OR uut_a_4_5 /= "000000001101011011100000011" OR uut_a_5_0 /= "111111111111011110001111101" OR uut_a_5_1 /= "000000001100101010001000101" OR uut_a_5_2 /= "000000000000010000111000001" OR uut_a_5_3 /= "111111111111011100001011111" OR uut_a_5_4 /= "000000001101011011100000011" OR uut_a_5_5 /= "000000000000010001111010000" THEN
              FAIL <= '1';
              FAIL_NUM <= "00001100";
              state <= "11111101";
            ELSE
              state <= "00011010";
            END IF;
            uut_rst <= '0';
          WHEN "00011010" =>
            uut_coord_shift <= "0110";
            uut_x <= "000001101001";
            uut_y <= "111110011011";
            uut_fx <= "0011111011";
            uut_fy <= "0011110010";
            uut_ft <= "0000111111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000101000100000000000" OR uut_a_0_1 /= "111110100010010110000000000" OR uut_a_0_2 /= "000000010100010000000000000" OR uut_a_0_3 /= "111111111101000000110000000" OR uut_a_0_4 /= "000000110111010010001000000" OR uut_a_0_5 /= "111111110100000011000000000" OR uut_a_1_0 /= "111111111101000100101100000" OR uut_a_1_1 /= "000000110110001001010010000" OR uut_a_1_2 /= "111111110100010010110000000" OR uut_a_1_3 /= "000000000001101110100100010" OR uut_a_1_4 /= "111111100000000010100001011" OR uut_a_1_5 /= "000000000110111010010001000" OR uut_a_2_0 /= "000000000000101000100000000" OR uut_a_2_1 /= "111111110100010010110000000" OR uut_a_2_2 /= "000000000010100010000000000" OR uut_a_2_3 /= "111111111111101000000110000" OR uut_a_2_4 /= "000000000110111010010001000" OR uut_a_2_5 /= "111111111110100000011000000" OR uut_a_3_0 /= "111111111101000000110000000" OR uut_a_3_1 /= "000000110111010010001000000" OR uut_a_3_2 /= "111111110100000011000000000" OR uut_a_3_3 /= "000000000001110000111001000" OR uut_a_3_4 /= "111111011111010111100001100" OR uut_a_3_5 /= "000000000111000011100100000" OR uut_a_4_0 /= "000000000001101110100100010" OR uut_a_4_1 /= "111111100000000010100001011" OR uut_a_4_2 /= "000000000110111010010001000" OR uut_a_4_3 /= "111111111110111110101111000" OR uut_a_4_4 /= "000000010010110111011001101" OR uut_a_4_5 /= "111111111011111010111100001" OR uut_a_5_0 /= "111111111111101000000110000" OR uut_a_5_1 /= "000000000110111010010001000" OR uut_a_5_2 /= "111111111110100000011000000" OR uut_a_5_3 /= "000000000000001110000111001" OR uut_a_5_4 /= "111111111011111010111100001" OR uut_a_5_5 /= "000000000000111000011100100" THEN
              FAIL <= '1';
              FAIL_NUM <= "00001101";
              state <= "11111101";
            ELSE
              state <= "00011011";
            END IF;
            uut_rst <= '0';
          WHEN "00011011" =>
            uut_coord_shift <= "0110";
            uut_x <= "111110110000";
            uut_y <= "000000011000";
            uut_fx <= "1100110011";
            uut_fy <= "1010001001";
            uut_ft <= "1011011010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000100111110110010000000" OR uut_a_0_1 /= "010001101111101010001000000" OR uut_a_0_2 /= "101111100000000010011000000" OR uut_a_0_3 /= "000000100100001100101100000" OR uut_a_0_4 /= "010000000111101001100110000" OR uut_a_0_5 /= "110001000000101111110010000" OR uut_a_1_0 /= "000000100011011111010100010" OR uut_a_1_1 /= "001111110011011100100001001" OR uut_a_1_2 /= "110001010011100010000111011" OR uut_a_1_3 /= "000000100000001111010011001" OR uut_a_1_4 /= "001110010110110100000010110" OR uut_a_1_5 /= "110010101001101010100011100" OR uut_a_2_0 /= "111111011111000000000100110" OR uut_a_2_1 /= "110001010011100010000111011" OR uut_a_2_2 /= "001101101010011110000010001" OR uut_a_2_3 /= "111111100010000001011111100" OR uut_a_2_4 /= "110010101001101010100011100" OR uut_a_2_5 /= "001100011010011000011011100" OR uut_a_3_0 /= "000000100100001100101100000" OR uut_a_3_1 /= "010000000111101001100110000" OR uut_a_3_2 /= "110001000000101111110010000" OR uut_a_3_3 /= "000000100000111000100001000" OR uut_a_3_4 /= "001110101001001010101100100" OR uut_a_3_5 /= "110010011000100110010101100" OR uut_a_4_0 /= "000000100000001111010011001" OR uut_a_4_1 /= "001110010110110100000010110" OR uut_a_4_2 /= "110010101001101010100011100" OR uut_a_4_3 /= "000000011101010010010101011" OR uut_a_4_4 /= "001101000010101010100001101" OR uut_a_4_5 /= "110011110111111010001001001" OR uut_a_5_0 /= "111111100010000001011111100" OR uut_a_5_1 /= "110010101001101010100011100" OR uut_a_5_2 /= "001100011010011000011011100" OR uut_a_5_3 /= "111111100100110001001100101" OR uut_a_5_4 /= "110011110111111010001001001" OR uut_a_5_5 /= "001011010001101000010000001" THEN
              FAIL <= '1';
              FAIL_NUM <= "00001110";
              state <= "11111101";
            ELSE
              state <= "00011100";
            END IF;
            uut_rst <= '0';
          WHEN "00011100" =>
            uut_coord_shift <= "0110";
            uut_x <= "000001100101";
            uut_y <= "111110010011";
            uut_fx <= "1011111000";
            uut_fy <= "1000110111";
            uut_ft <= "1111000100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000110011011011111001000" OR uut_a_0_1 /= "000110000001110001001011100" OR uut_a_0_2 /= "000011100111011101100000100" OR uut_a_0_3 /= "111111001110011110000010000" OR uut_a_0_4 /= "111010001100100001001111000" OR uut_a_0_5 /= "111100100001000111001001000" OR uut_a_1_0 /= "000000001100000011100010010" OR uut_a_1_1 /= "000001011010011010100001101" OR uut_a_1_2 /= "000000110110001111111010100" OR uut_a_1_3 /= "111111110100011001000010011" OR uut_a_1_4 /= "111110101000111011110010100" OR uut_a_1_5 /= "111111001011110000101011000" OR uut_a_2_0 /= "000000000111001110111011000" OR uut_a_2_1 /= "000000110110001111111010100" OR uut_a_2_2 /= "000000100000100011001001100" OR uut_a_2_3 /= "111111111001000010001110010" OR uut_a_2_4 /= "111111001011110000101011000" OR uut_a_2_5 /= "111111100000101010000000010" OR uut_a_3_0 /= "111111001110011110000010000" OR uut_a_3_1 /= "111010001100100001001111000" OR uut_a_3_2 /= "111100100001000111001001000" OR uut_a_3_3 /= "000000101111101100100100000" OR uut_a_3_4 /= "000101100101101110001110000" OR uut_a_3_5 /= "000011010110101000100010000" OR uut_a_4_0 /= "111111110100011001000010011" OR uut_a_4_1 /= "111110101000111011110010100" OR uut_a_4_2 /= "111111001011110000101011000" OR uut_a_4_3 /= "000000001011001011011100011" OR uut_a_4_4 /= "000001010011110101110101010" OR uut_a_4_5 /= "000000110010010011011111111" OR uut_a_5_0 /= "111111111001000010001110010" OR uut_a_5_1 /= "111111001011110000101011000" OR uut_a_5_2 /= "111111100000101010000000010" OR uut_a_5_3 /= "000000000110101101010001000" OR uut_a_5_4 /= "000000110010010011011111111" OR uut_a_5_5 /= "000000011110001011101100110" THEN
              FAIL <= '1';
              FAIL_NUM <= "00001111";
              state <= "11111101";
            ELSE
              state <= "00011101";
            END IF;
            uut_rst <= '0';
          WHEN "00011101" =>
            uut_coord_shift <= "0110";
            uut_x <= "111110000100";
            uut_y <= "000001100101";
            uut_fx <= "1011001001";
            uut_fy <= "1001100000";
            uut_ft <= "1100111011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000100001001111100001000" OR uut_a_0_1 /= "000111110010101000101111000" OR uut_a_0_2 /= "110001101101110101010100100" OR uut_a_0_3 /= "000000101000000101101101000" OR uut_a_0_4 /= "001001011001010101100011000" OR uut_a_0_5 /= "101110110001100011001010100" OR uut_a_1_0 /= "000000001111100101010001011" OR uut_a_1_1 /= "000011101001101111000110000" OR uut_a_1_2 /= "111001010011011110111111100" OR uut_a_1_3 /= "000000010010110010101011000" OR uut_a_1_4 /= "000100011001111000000110011" OR uut_a_1_5 /= "110111111011001110011110111" OR uut_a_2_0 /= "111111100011011011101010101" OR uut_a_2_1 /= "111001010011011110111111100" OR uut_a_2_2 /= "001100010001100111001011011" OR uut_a_2_3 /= "111111011101100011000110010" OR uut_a_2_4 /= "110111111011001110011110111" OR uut_a_2_5 /= "001110110011011010110001111" OR uut_a_3_0 /= "000000101000000101101101000" OR uut_a_3_1 /= "001001011001010101100011000" OR uut_a_3_2 /= "101110110001100011001010100" OR uut_a_3_3 /= "000000110000010110001001000" OR uut_a_3_4 /= "001011010101001100000111000" OR uut_a_3_5 /= "101011001110011111001000100" OR uut_a_4_0 /= "000000010010110010101011000" OR uut_a_4_1 /= "000100011001111000000110011" OR uut_a_4_2 /= "110111111011001110011110111" OR uut_a_4_3 /= "000000010110101010011000001" OR uut_a_4_4 /= "000101010011111011101011010" OR uut_a_4_5 /= "110110010000110010100101111" OR uut_a_5_0 /= "111111011101100011000110010" OR uut_a_5_1 /= "110111111011001110011110111" OR uut_a_5_2 /= "001110110011011010110001111" OR uut_a_5_3 /= "111111010110011100111110010" OR uut_a_5_4 /= "110110010000110010100101111" OR uut_a_5_5 /= "010001110110100011001111101" THEN
              FAIL <= '1';
              FAIL_NUM <= "00010000";
              state <= "11111101";
            ELSE
              state <= "00011110";
            END IF;
            uut_rst <= '0';
          WHEN "00011110" =>
            uut_coord_shift <= "0110";
            uut_x <= "111111110101";
            uut_y <= "111110011011";
            uut_fx <= "0111111011";
            uut_fy <= "1101010100";
            uut_ft <= "1100110000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000011000100000" OR uut_a_0_1 /= "000000000001000100111010000" OR uut_a_0_2 /= "000000000000110111001000000" OR uut_a_0_3 /= "111111111110110111110100000" OR uut_a_0_4 /= "111111100110100111110010000" OR uut_a_0_5 /= "111111101011101100101000000" OR uut_a_1_0 /= "000000000000000010001001110" OR uut_a_1_1 /= "000000000000110000011100110" OR uut_a_1_2 /= "000000000000100110110000101" OR uut_a_1_3 /= "111111111111001101001111100" OR uut_a_1_4 /= "111111101110001001111110001" OR uut_a_1_5 /= "111111110001101110011000001" OR uut_a_2_0 /= "000000000000000001101110010" OR uut_a_2_1 /= "000000000000100110110000101" OR uut_a_2_2 /= "000000000000011111000000100" OR uut_a_2_3 /= "111111111111010111011001010" OR uut_a_2_4 /= "111111110001101110011000001" OR uut_a_2_5 /= "111111110100100101000110100" OR uut_a_3_0 /= "111111111110110111110100000" OR uut_a_3_1 /= "111111100110100111110010000" OR uut_a_3_2 /= "111111101011101100101000000" OR uut_a_3_3 /= "000000011010100101100100000" OR uut_a_3_4 /= "001001010110001101001010000" OR uut_a_3_5 /= "000111011110100100001000000" OR uut_a_4_0 /= "111111111111001101001111100" OR uut_a_4_1 /= "111111101110001001111110001" OR uut_a_4_2 /= "111111110001101110011000001" OR uut_a_4_3 /= "000000010010101100011010010" OR uut_a_4_4 /= "000110100100100111010000000" OR uut_a_4_5 /= "000101010000011111011001101" OR uut_a_5_0 /= "111111111111010111011001010" OR uut_a_5_1 /= "111111110001101110011000001" OR uut_a_5_2 /= "111111110100100101000110100" OR uut_a_5_3 /= "000000001110111101001000010" OR uut_a_5_4 /= "000101010000011111011001101" OR uut_a_5_5 /= "000100001101001100010100100" THEN
              FAIL <= '1';
              FAIL_NUM <= "00010001";
              state <= "11111101";
            ELSE
              state <= "00011111";
            END IF;
            uut_rst <= '0';
          WHEN "00011111" =>
            uut_coord_shift <= "0110";
            uut_x <= "111110010000";
            uut_y <= "111111001101";
            uut_fx <= "1000101111";
            uut_fy <= "0000000110";
            uut_ft <= "0100001100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000110001011100000100000" OR uut_a_0_1 /= "101110001110111010100100000" OR uut_a_0_2 /= "101000110100110110001000000" OR uut_a_0_3 /= "111111101001101100101010000" OR uut_a_0_4 /= "001000000000111100111010000" OR uut_a_0_5 /= "001010011101000100010100000" OR uut_a_1_0 /= "111111011100011101110101001" OR uut_a_1_1 /= "001100110001010001111010001" OR uut_a_1_2 /= "010000101010000001000110010" OR uut_a_1_3 /= "000000010000000001111001110" OR uut_a_1_4 /= "111010001111010100001110010" OR uut_a_1_5 /= "111000011111000110111001101" OR uut_a_2_0 /= "111111010001101001101100010" OR uut_a_2_1 /= "010000101010000001000110010" OR uut_a_2_2 /= "010101101110011101010000100" OR uut_a_2_3 /= "000000010100111010001000101" OR uut_a_2_4 /= "111000011111000110111001101" OR uut_a_2_5 /= "110110001100101111111101010" OR uut_a_3_0 /= "111111101001101100101010000" OR uut_a_3_1 /= "001000000000111100111010000" OR uut_a_3_2 /= "001010011101000100010100000" OR uut_a_3_3 /= "000000001010000011111001000" OR uut_a_3_4 /= "111100011000100110100001000" OR uut_a_3_5 /= "111011010010001011010010000" OR uut_a_4_0 /= "000000010000000001111001110" OR uut_a_4_1 /= "111010001111010100001110010" OR uut_a_4_2 /= "111000011111000110111001101" OR uut_a_4_3 /= "111111111000110001001101000" OR uut_a_4_4 /= "000010100110010100010100010" OR uut_a_4_5 /= "000011011000111011111001000" OR uut_a_5_0 /= "000000010100111010001000101" OR uut_a_5_1 /= "111000011111000110111001101" OR uut_a_5_2 /= "110110001100101111111101010" OR uut_a_5_3 /= "111111110110100100010110100" OR uut_a_5_4 /= "000011011000111011111001000" OR uut_a_5_5 /= "000100011010111101011011001" THEN
              FAIL <= '1';
              FAIL_NUM <= "00010010";
              state <= "11111101";
            ELSE
              state <= "00100000";
            END IF;
            uut_rst <= '0';
          WHEN "00100000" =>
            uut_coord_shift <= "0110";
            uut_x <= "000000100001";
            uut_y <= "111110011000";
            uut_fx <= "1001010011";
            uut_fy <= "0100011100";
            uut_ft <= "0110011111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000101101001000000000" OR uut_a_0_1 /= "111111000100110001100000000" OR uut_a_0_2 /= "111111110100101110000000000" OR uut_a_0_3 /= "111111101101111101110000000" OR uut_a_0_4 /= "000010111101010111101000000" OR uut_a_0_5 /= "000000100100000100100000000" OR uut_a_1_0 /= "111111111110001001100011000" OR uut_a_1_1 /= "000000010011011011110000100" OR uut_a_1_2 /= "000000000011101100111010000" OR uut_a_1_3 /= "000000000101111010101111010" OR uut_a_1_4 /= "111111000001110111001111111" OR uut_a_1_5 /= "111111110100001010100001100" OR uut_a_2_0 /= "111111111111101001011100000" OR uut_a_2_1 /= "000000000011101100111010000" OR uut_a_2_2 /= "000000000000101101001000000" OR uut_a_2_3 /= "000000000001001000001001000" OR uut_a_2_4 /= "111111110100001010100001100" OR uut_a_2_5 /= "111111111101101111101110000" OR uut_a_3_0 /= "111111101101111101110000000" OR uut_a_3_1 /= "000010111101010111101000000" OR uut_a_3_2 /= "000000100100000100100000000" OR uut_a_3_3 /= "000000111001101010100100000" OR uut_a_3_4 /= "110110100010100001000110000" OR uut_a_3_5 /= "111110001100101010111000000" OR uut_a_4_0 /= "000000000101111010101111010" OR uut_a_4_1 /= "111111000001110111001111111" OR uut_a_4_2 /= "111111110100001010100001100" OR uut_a_4_3 /= "111111101101000101000010001" OR uut_a_4_4 /= "000011000110101011001001000" OR uut_a_4_5 /= "000000100101110101111011101" OR uut_a_5_0 /= "000000000001001000001001000" OR uut_a_5_1 /= "111111110100001010100001100" OR uut_a_5_2 /= "111111111101101111101110000" OR uut_a_5_3 /= "111111111100011001010101110" OR uut_a_5_4 /= "000000100101110101111011101" OR uut_a_5_5 /= "000000000111001101010100100" THEN
              FAIL <= '1';
              FAIL_NUM <= "00010011";
              state <= "11111101";
            ELSE
              state <= "00100001";
            END IF;
            uut_rst <= '0';
          WHEN "00100001" =>
            uut_coord_shift <= "0110";
            uut_x <= "000000001000";
            uut_y <= "111110011100";
            uut_fx <= "0101001110";
            uut_fy <= "1101011010";
            uut_ft <= "1100101101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000010111110001000000" OR uut_a_0_1 /= "000000010110010001111100000" OR uut_a_0_2 /= "000010000101101011101000000" OR uut_a_0_3 /= "000000000001000011000010000" OR uut_a_0_4 /= "000000000111110110101111000" OR uut_a_0_5 /= "000000101111001000011010000" OR uut_a_1_0 /= "000000000000010110010001111" OR uut_a_1_1 /= "000000000010100111000110100" OR uut_a_1_2 /= "000000001111101010100111001" OR uut_a_1_3 /= "000000000000000111110110101" OR uut_a_1_4 /= "000000000000111010111010100" OR uut_a_1_5 /= "000000000101100001011111000" OR uut_a_2_0 /= "000000000010000101101011101" OR uut_a_2_1 /= "000000001111101010100111001" OR uut_a_2_2 /= "000001011101111111101011001" OR uut_a_2_3 /= "000000000000101111001000011" OR uut_a_2_4 /= "000000000101100001011111000" OR uut_a_2_5 /= "000000100001001000111010010" OR uut_a_3_0 /= "000000000001000011000010000" OR uut_a_3_1 /= "000000000111110110101111000" OR uut_a_3_2 /= "000000101111001000011010000" OR uut_a_3_3 /= "000000000000010111101000100" OR uut_a_3_4 /= "000000000010110001001111110" OR uut_a_3_5 /= "000000010000100111011110100" OR uut_a_4_0 /= "000000000000000111110110101" OR uut_a_4_1 /= "000000000000111010111010100" OR uut_a_4_2 /= "000000000101100001011111000" OR uut_a_4_3 /= "000000000000000010110001001" OR uut_a_4_4 /= "000000000000010100110001010" OR uut_a_4_5 /= "000000000001111100101000000" OR uut_a_5_0 /= "000000000000101111001000011" OR uut_a_5_1 /= "000000000101100001011111000" OR uut_a_5_2 /= "000000100001001000111010010" OR uut_a_5_3 /= "000000000000010000100111011" OR uut_a_5_4 /= "000000000001111100101000000" OR uut_a_5_5 /= "000000001011101011110000011" THEN
              FAIL <= '1';
              FAIL_NUM <= "00010100";
              state <= "11111101";
            ELSE
              state <= "00100010";
            END IF;
            uut_rst <= '0';
          WHEN "00100010" =>
            uut_coord_shift <= "0110";
            uut_x <= "000000111111";
            uut_y <= "111110000011";
            uut_fx <= "1000110010";
            uut_fy <= "0010101100";
            uut_ft <= "0001101010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000011101001110100100" OR uut_a_0_1 /= "111101101010001101010111100" OR uut_a_0_2 /= "000001001010111001010100010" OR uut_a_0_3 /= "111111110111011000100100000" OR uut_a_0_4 /= "000101100001010000111100000" OR uut_a_0_5 /= "111101001111010111100010000" OR uut_a_1_0 /= "111111111101101010001101010" OR uut_a_1_1 /= "000001011111111101011011111" OR uut_a_1_2 /= "111111010000000001010010000" OR uut_a_1_3 /= "000000000101100001010000111" OR uut_a_1_4 /= "111100011101101100001001100" OR uut_a_1_5 /= "000001110001001001111011001" OR uut_a_2_0 /= "000000000001001010111001010" OR uut_a_2_1 /= "111111010000000001010010000" OR uut_a_2_2 /= "000000010111111111010110111" OR uut_a_2_3 /= "111111111101001111010111100" OR uut_a_2_4 /= "000001110001001001111011001" OR uut_a_2_5 /= "111111000111011011000010011" OR uut_a_3_0 /= "111111110111011000100100000" OR uut_a_3_1 /= "000101100001010000111100000" OR uut_a_3_2 /= "111101001111010111100010000" OR uut_a_3_3 /= "000000010100010100100000000" OR uut_a_3_4 /= "110010111110110111100000000" OR uut_a_3_5 /= "000110100000100100010000000" OR uut_a_4_0 /= "000000000101100001010000111" OR uut_a_4_1 /= "111100011101101100001001100" OR uut_a_4_2 /= "000001110001001001111011001" OR uut_a_4_3 /= "111111110010111110110111100" OR uut_a_4_4 /= "001000010101101110011100100" OR uut_a_4_5 /= "111011110101001000110001110" OR uut_a_5_0 /= "111111111101001111010111100" OR uut_a_5_1 /= "000001110001001001111011001" OR uut_a_5_2 /= "111111000111011011000010011" OR uut_a_5_3 /= "000000000110100000100100010" OR uut_a_5_4 /= "111011110101001000110001110" OR uut_a_5_5 /= "000010000101011011100111001" THEN
              FAIL <= '1';
              FAIL_NUM <= "00010101";
              state <= "11111101";
            ELSE
              state <= "00100011";
            END IF;
            uut_rst <= '0';
          WHEN "00100011" =>
            uut_coord_shift <= "0110";
            uut_x <= "000000000110";
            uut_y <= "000000111010";
            uut_fx <= "0011010100";
            uut_fy <= "0100100000";
            uut_ft <= "1100100111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000101011111001000000" OR uut_a_0_1 /= "000101010110111001010100000" OR uut_a_0_2 /= "000000011011011011101000000" OR uut_a_0_3 /= "000000001101001110010110000" OR uut_a_0_4 /= "001100111010100000011111000" OR uut_a_0_5 /= "000001000010000111101110000" OR uut_a_1_0 /= "000000000101010110111001010" OR uut_a_1_1 /= "000101001110110110111110000" OR uut_a_1_2 /= "000000011010110010011110100" OR uut_a_1_3 /= "000000001100111010100000011" OR uut_a_1_4 /= "001100100111001000101110010" OR uut_a_1_5 /= "000001000000100100100010011" OR uut_a_2_0 /= "000000000000011011011011101" OR uut_a_2_1 /= "000000011010110010011110100" OR uut_a_2_2 /= "000000000010001001001010001" OR uut_a_2_3 /= "000000000001000010000111101" OR uut_a_2_4 /= "000001000000100100100010011" OR uut_a_2_5 /= "000000000101001010100110100" OR uut_a_3_0 /= "000000001101001110010110000" OR uut_a_3_1 /= "001100111010100000011111000" OR uut_a_3_2 /= "000001000010000111101110000" OR uut_a_3_3 /= "000000011111111000000000100" OR uut_a_3_4 /= "011111001000001100011111010" OR uut_a_3_5 /= "000010011111011000000010100" OR uut_a_4_0 /= "000000001100111010100000011" OR uut_a_4_1 /= "001100100111001000101110010" OR uut_a_4_2 /= "000001000000100100100010011" OR uut_a_4_3 /= "000000011111001000001100011" OR uut_a_4_4 /= "011110011001100000001100100" OR uut_a_4_5 /= "000010011011101000111110011" OR uut_a_5_0 /= "000000000001000010000111101" OR uut_a_5_1 /= "000001000000100100100010011" OR uut_a_5_2 /= "000000000101001010100110100" OR uut_a_5_3 /= "000000000010011111011000000" OR uut_a_5_4 /= "000010011011101000111110011" OR uut_a_5_5 /= "000000001100011100111000001" THEN
              FAIL <= '1';
              FAIL_NUM <= "00010110";
              state <= "11111101";
            ELSE
              state <= "00100100";
            END IF;
            uut_rst <= '0';
          WHEN "00100100" =>
            uut_coord_shift <= "0110";
            uut_x <= "000000110001";
            uut_y <= "000000001110";
            uut_fx <= "1110010110";
            uut_fy <= "1000111111";
            uut_ft <= "0100011111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000001000111001100010000" OR uut_a_0_1 /= "111110100010100011111011000" OR uut_a_0_2 /= "111111010111111101000111000" OR uut_a_0_3 /= "000000001010101111101010000" OR uut_a_0_4 /= "111110001111001011100111000" OR uut_a_0_5 /= "111111001111101001100011000" OR uut_a_1_0 /= "111111111110100010100011111" OR uut_a_1_1 /= "000000001111010101000110110" OR uut_a_1_2 /= "000000000110100100011110010" OR uut_a_1_3 /= "111111111110001111001011100" OR uut_a_1_4 /= "000000010010100000100110000" OR uut_a_1_5 /= "000000000111111011101011110" OR uut_a_2_0 /= "111111111111010111111101000" OR uut_a_2_1 /= "000000000110100100011110010" OR uut_a_2_2 /= "000000000010110100001101000" OR uut_a_2_3 /= "111111111111001111101001100" OR uut_a_2_4 /= "000000000111111011101011110" OR uut_a_2_5 /= "000000000011011001100101000" OR uut_a_3_0 /= "000000001010101111101010000" OR uut_a_3_1 /= "111110001111001011100111000" OR uut_a_3_2 /= "111111001111101001100011000" OR uut_a_3_3 /= "000000001100111110010010000" OR uut_a_3_4 /= "111101110111110010000011000" OR uut_a_3_5 /= "111111000101100111101111000" OR uut_a_4_0 /= "111111111110001111001011100" OR uut_a_4_1 /= "000000010010100000100110000" OR uut_a_4_2 /= "000000000111111011101011110" OR uut_a_4_3 /= "111111111101110111110010000" OR uut_a_4_4 /= "000000010110010110010010100" OR uut_a_4_5 /= "000000001001100100111110110" OR uut_a_5_0 /= "111111111111001111101001100" OR uut_a_5_1 /= "000000000111111011101011110" OR uut_a_5_2 /= "000000000011011001100101000" OR uut_a_5_3 /= "111111111111000101100111101" OR uut_a_5_4 /= "000000001001100100111110110" OR uut_a_5_5 /= "000000000100000110101101001" THEN
              FAIL <= '1';
              FAIL_NUM <= "00010111";
              state <= "11111101";
            ELSE
              state <= "00100101";
            END IF;
            uut_rst <= '0';
          WHEN "00100101" =>
            uut_coord_shift <= "0110";
            uut_x <= "111111010111";
            uut_y <= "000000011011";
            uut_fx <= "0011110111";
            uut_fy <= "1001101011";
            uut_ft <= "1010000011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000011001001010010010000" OR uut_a_0_1 /= "101111111000011010011110000" OR uut_a_0_2 /= "111001000111101100000101000" OR uut_a_0_3 /= "111111111110110001111110000" OR uut_a_0_4 /= "000000110001111111010010000" OR uut_a_0_5 /= "000000010101010101100011000" OR uut_a_1_0 /= "111111101111111000011010011" OR uut_a_1_1 /= "001010010100110111000010110" OR uut_a_1_2 /= "000100011010000100110000110" OR uut_a_1_3 /= "000000000000110001111111010" OR uut_a_1_4 /= "111111011111111110011101011" OR uut_a_1_5 /= "111111110010010101001100100" OR uut_a_2_0 /= "111111111001000111101100000" OR uut_a_2_1 /= "000100011010000100110000110" OR uut_a_2_2 /= "000001111000011001011100101" OR uut_a_2_3 /= "000000000000010101010101100" OR uut_a_2_4 /= "111111110010010101001100100" OR uut_a_2_5 /= "111111111010001010100110111" OR uut_a_3_0 /= "111111111110110001111110000" OR uut_a_3_1 /= "000000110001111111010010000" OR uut_a_3_2 /= "000000010101010101100011000" OR uut_a_3_3 /= "000000000000000011110010000" OR uut_a_3_4 /= "111111111101100100111110000" OR uut_a_3_5 /= "111111111110111101110101000" OR uut_a_4_0 /= "000000000000110001111111010" OR uut_a_4_1 /= "111111011111111110011101011" OR uut_a_4_2 /= "111111110010010101001100100" OR uut_a_4_3 /= "111111111111111101100100111" OR uut_a_4_4 /= "000000000001100011010100010" OR uut_a_4_5 /= "000000000000101010011001000" OR uut_a_5_0 /= "000000000000010101010101100" OR uut_a_5_1 /= "111111110010010101001100100" OR uut_a_5_2 /= "111111111010001010100110111" OR uut_a_5_3 /= "111111111111111110111101110" OR uut_a_5_4 /= "000000000000101010011001000" OR uut_a_5_5 /= "000000000000010010000110000" THEN
              FAIL <= '1';
              FAIL_NUM <= "00011000";
              state <= "11111101";
            ELSE
              state <= "00100110";
            END IF;
            uut_rst <= '0';
          WHEN "00100110" =>
            uut_coord_shift <= "0110";
            uut_x <= "000000001100";
            uut_y <= "111111111101";
            uut_fx <= "0110010000";
            uut_fy <= "0100110010";
            uut_ft <= "0011110000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000010101000001100000100" OR uut_a_0_1 /= "110010010111100001011011010" OR uut_a_0_2 /= "110011110110001000001101100" OR uut_a_0_3 /= "000000001001000111100110000" OR uut_a_0_4 /= "111010000101100100110111000" OR uut_a_0_5 /= "111010101110100111000010000" OR uut_a_1_0 /= "111111110010010111100001011" OR uut_a_1_1 /= "001000110101101111110100110" OR uut_a_1_2 /= "000111111000011001101011001" OR uut_a_1_3 /= "111111111010000101100100110" OR uut_a_1_4 /= "000011110101011000100110010" OR uut_a_1_5 /= "000011011010110001101100001" OR uut_a_2_0 /= "111111110011110110001000001" OR uut_a_2_1 /= "000111111000011001101011001" OR uut_a_2_2 /= "000111000001101101010000001" OR uut_a_2_3 /= "111111111010101110100111000" OR uut_a_2_4 /= "000011011010110001101100001" OR uut_a_2_5 /= "000011000011000011011011110" OR uut_a_3_0 /= "000000001001000111100110000" OR uut_a_3_1 /= "111010000101100100110111000" OR uut_a_3_2 /= "111010101110100111000010000" OR uut_a_3_3 /= "000000000011111101001000000" OR uut_a_3_4 /= "111101011011110111010100000" OR uut_a_3_5 /= "111101101101101010011000000" OR uut_a_4_0 /= "111111111010000101100100110" OR uut_a_4_1 /= "000011110101011000100110010" OR uut_a_4_2 /= "000011011010110001101100001" OR uut_a_4_3 /= "111111111101011011110111010" OR uut_a_4_4 /= "000001101010011011101000100" OR uut_a_4_5 /= "000001011110111001000001011" OR uut_a_5_0 /= "111111111010101110100111000" OR uut_a_5_1 /= "000011011010110001101100001" OR uut_a_5_2 /= "000011000011000011011011110" OR uut_a_5_3 /= "111111111101101101101010011" OR uut_a_5_4 /= "000001011110111001000001011" OR uut_a_5_5 /= "000001010100100110100000001" THEN
              FAIL <= '1';
              FAIL_NUM <= "00011001";
              state <= "11111101";
            ELSE
              state <= "00100111";
            END IF;
            uut_rst <= '0';
          WHEN "00100111" =>
            uut_coord_shift <= "0110";
            uut_x <= "111110001110";
            uut_y <= "111110010011";
            uut_fx <= "1001011011";
            uut_fy <= "0100110010";
            uut_ft <= "0111000110";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000111101100001100100" OR uut_a_0_1 /= "000110010011110000010000010" OR uut_a_0_2 /= "111001111011101000001000110" OR uut_a_0_3 /= "000000000111011010100011000" OR uut_a_0_4 /= "000110000101010001101101100" OR uut_a_0_5 /= "111010001001100011011000100" OR uut_a_1_0 /= "000000000110010011110000010" OR uut_a_1_1 /= "000101001011001101000101010" OR uut_a_1_2 /= "111011000001011010011011001" OR uut_a_1_3 /= "000000000110000101010001101" OR uut_a_1_4 /= "000100111111010101000001110" OR uut_a_1_5 /= "111011001100110101100001100" OR uut_a_2_0 /= "111111111001111011101000001" OR uut_a_2_1 /= "111011000001011010011011001" OR uut_a_2_2 /= "000100110010011100110101000" OR uut_a_2_3 /= "111111111010001001100011011" OR uut_a_2_4 /= "111011001100110101100001100" OR uut_a_2_5 /= "000100100111011101100101001" OR uut_a_3_0 /= "000000000111011010100011000" OR uut_a_3_1 /= "000110000101010001101101100" OR uut_a_3_2 /= "111010001001100011011000100" OR uut_a_3_3 /= "000000000111001001100010000" OR uut_a_3_4 /= "000101110111010100011001000" OR uut_a_3_5 /= "111010010110111110101011000" OR uut_a_4_0 /= "000000000110000101010001101" OR uut_a_4_1 /= "000100111111010101000001110" OR uut_a_4_2 /= "111011001100110101100001100" OR uut_a_4_3 /= "000000000101110111010100011" OR uut_a_4_4 /= "000100110011111000001110100" OR uut_a_4_5 /= "111011010111110110011010010" OR uut_a_5_0 /= "111111111010001001100011011" OR uut_a_5_1 /= "111011001100110101100001100" OR uut_a_5_2 /= "000100100111011101100101001" OR uut_a_5_3 /= "111111111010010110111110101" OR uut_a_5_4 /= "111011010111110110011010010" OR uut_a_5_5 /= "000100011100110111100011000" THEN
              FAIL <= '1';
              FAIL_NUM <= "00011010";
              state <= "11111101";
            ELSE
              state <= "00101000";
            END IF;
            uut_rst <= '0';
          WHEN "00101000" =>
            uut_coord_shift <= "0111";
            uut_x <= "000001011110";
            uut_y <= "111101000100";
            uut_fx <= "0011100100";
            uut_fy <= "1001110001";
            uut_ft <= "1001111000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000101001000010100100" OR uut_a_0_1 /= "111100110010110011001100000" OR uut_a_0_2 /= "000000111101100011110110000" OR uut_a_0_3 /= "000000001001011000100101100" OR uut_a_0_4 /= "111010001000101000100100000" OR uut_a_0_5 /= "000001110000100111000010000" OR uut_a_1_0 /= "111111111100110010110011001" OR uut_a_1_1 /= "000010000000010000000000100" OR uut_a_1_2 /= "111111011001100001100110010" OR uut_a_1_3 /= "111111111010001000101000100" OR uut_a_1_4 /= "000011101010100110101001100" OR uut_a_1_5 /= "111110111001100111100110110" OR uut_a_2_0 /= "000000000000111101100011110" OR uut_a_2_1 /= "111111011001100001100110010" OR uut_a_2_2 /= "000000001011100010101110001" OR uut_a_2_3 /= "000000000001110000100111000" OR uut_a_2_4 /= "111110111001100111100110110" OR uut_a_2_5 /= "000000010101000111010100011" OR uut_a_3_0 /= "000000001001011000100101100" OR uut_a_3_1 /= "111010001000101000100100000" OR uut_a_3_2 /= "000001110000100111000010000" OR uut_a_3_3 /= "000000010001001010101000100" OR uut_a_3_4 /= "110101010001010110101100000" OR uut_a_3_5 /= "000011001101111111100110000" OR uut_a_4_0 /= "111111111010001000101000100" OR uut_a_4_1 /= "000011101010100110101001100" OR uut_a_4_2 /= "111110111001100111100110110" OR uut_a_4_3 /= "111111110101010001010110101" OR uut_a_4_4 /= "000110101101001001110100100" OR uut_a_4_5 /= "111101111111010000010000010" OR uut_a_5_0 /= "000000000001110000100111000" OR uut_a_5_1 /= "111110111001100111100110110" OR uut_a_5_2 /= "000000010101000111010100011" OR uut_a_5_3 /= "000000000011001101111111100" OR uut_a_5_4 /= "111101111111010000010000010" OR uut_a_5_5 /= "000000100110100111111011001" THEN
              FAIL <= '1';
              FAIL_NUM <= "00011011";
              state <= "11111101";
            ELSE
              state <= "00101001";
            END IF;
            uut_rst <= '0';
          WHEN "00101001" =>
            uut_coord_shift <= "0111";
            uut_x <= "000001001000";
            uut_y <= "111110101001";
            uut_fx <= "0010011110";
            uut_fy <= "0011111111";
            uut_ft <= "0001010101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000001000100000100000000" OR uut_a_0_1 /= "000110101101101001010000000" OR uut_a_0_2 /= "111000110000010100110000000" OR uut_a_0_3 /= "000000001110101110100100000" OR uut_a_0_4 /= "001011100111101111011010000" OR uut_a_0_5 /= "110011011101010110010110000" OR uut_a_1_0 /= "000000000110101101101001010" OR uut_a_1_1 /= "000101010011000001000011001" OR uut_a_1_2 /= "111010010010001000010111111" OR uut_a_1_3 /= "000000001011100111101111011" OR uut_a_1_4 /= "001001001010110110111010000" OR uut_a_1_5 /= "110110000110101010001000010" OR uut_a_2_0 /= "111111111000110000010100110" OR uut_a_2_1 /= "111010010010001000010111111" OR uut_a_2_2 /= "000110001010110110010101001" OR uut_a_2_3 /= "111111110011011101010110010" OR uut_a_2_4 /= "110110000110101010001000010" OR uut_a_2_5 /= "001010101011100000011110010" OR uut_a_3_0 /= "000000001110101110100100000" OR uut_a_3_1 /= "001011100111101111011010000" OR uut_a_3_2 /= "110011011101010110010110000" OR uut_a_3_3 /= "000000011001011111101000100" OR uut_a_3_4 /= "010100000111011101011101010" OR uut_a_3_5 /= "101010010010100100000000110" OR uut_a_4_0 /= "000000001011100111101111011" OR uut_a_4_1 /= "001001001010110110111010000" OR uut_a_4_2 /= "110110000110101010001000010" OR uut_a_4_3 /= "000000010100000111011101011" OR uut_a_4_4 /= "001111110111111000101111100" OR uut_a_4_5 /= "101110110111101001011010100" OR uut_a_5_0 /= "111111110011011101010110010" OR uut_a_5_1 /= "110110000110101010001000010" OR uut_a_5_2 /= "001010101011100000011110010" OR uut_a_5_3 /= "111111101010010010100100000" OR uut_a_5_4 /= "101110110111101001011010100" OR uut_a_5_5 /= "010010011111001100010101010" THEN
              FAIL <= '1';
              FAIL_NUM <= "00011100";
              state <= "11111101";
            ELSE
              state <= "00101010";
            END IF;
            uut_rst <= '0';
          WHEN "00101010" =>
            uut_coord_shift <= "0111";
            uut_x <= "000001111010";
            uut_y <= "111101111001";
            uut_fx <= "0011110001";
            uut_fy <= "0111100010";
            uut_ft <= "0101111000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000001011110011101000100" OR uut_a_0_1 /= "110100100011111110110001000" OR uut_a_0_2 /= "001001010100001111011101010" OR uut_a_0_3 /= "000000001111110010110000000" OR uut_a_0_4 /= "110000101100110101100000000" OR uut_a_0_5 /= "001100011101100010111000000" OR uut_a_1_0 /= "111111110100100011111110110" OR uut_a_1_1 /= "001011000101001001001100100" OR uut_a_1_2 /= "110110111110011001000001101" OR uut_a_1_3 /= "111111110000101100110101100" OR uut_a_1_4 /= "001110110100100100001011000" OR uut_a_1_5 /= "110011111011011000001101110" OR uut_a_2_0 /= "000000001001010100001111011" OR uut_a_2_1 /= "110110111110011001000001101" OR uut_a_2_2 /= "000111010110011110001100100" OR uut_a_2_3 /= "000000001100011101100010111" OR uut_a_2_4 /= "110011111011011000001101110" OR uut_a_2_5 /= "001001110101010100000001001" OR uut_a_3_0 /= "000000001111110010110000000" OR uut_a_3_1 /= "110000101100110101100000000" OR uut_a_3_2 /= "001100011101100010111000000" OR uut_a_3_3 /= "000000010101001000000000000" OR uut_a_3_4 /= "101011100010010000000000000" OR uut_a_3_5 /= "010000101010110100000000000" OR uut_a_4_0 /= "111111110000101100110101100" OR uut_a_4_1 /= "001110110100100100001011000" OR uut_a_4_2 /= "110011111011011000001101110" OR uut_a_4_3 /= "111111101011100010010000000" OR uut_a_4_4 /= "010011110100110100100000000" OR uut_a_4_5 /= "101111110110100001101000000" OR uut_a_5_0 /= "000000001100011101100010111" OR uut_a_5_1 /= "110011111011011000001101110" OR uut_a_5_2 /= "001001110101010100000001001" OR uut_a_5_3 /= "000000010000101010110100000" OR uut_a_5_4 /= "101111110110100001101000000" OR uut_a_5_5 /= "001101001001110010000010000" THEN
              FAIL <= '1';
              FAIL_NUM <= "00011101";
              state <= "11111101";
            ELSE
              state <= "00101011";
            END IF;
            uut_rst <= '0';
          WHEN "00101011" =>
            uut_coord_shift <= "0111";
            uut_x <= "111100101101";
            uut_y <= "111110111100";
            uut_fx <= "1101111010";
            uut_fy <= "0010111101";
            uut_ft <= "0001100100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000011111011000001100100" OR uut_a_0_1 /= "111101010011011010111011010" OR uut_a_0_2 /= "100111001111011010001000110" OR uut_a_0_3 /= "111111110101010110101110000" OR uut_a_0_4 /= "000000111010100011000011000" OR uut_a_0_5 /= "001000011001100100101101000" OR uut_a_1_0 /= "111111111101010011011010111" OR uut_a_1_1 /= "000000001110110101001011111" OR uut_a_1_2 /= "000010001000001011010000001" OR uut_a_1_3 /= "000000000000111010100011000" OR uut_a_1_4 /= "111111111010111101111111001" OR uut_a_1_5 /= "111111010001110011010110001" OR uut_a_2_0 /= "111111100111001111011010001" OR uut_a_2_1 /= "000010001000001011010000001" OR uut_a_2_2 /= "010011100010010101111000000" OR uut_a_2_3 /= "000000001000011001100100101" OR uut_a_2_4 /= "111111010001110011010110001" OR uut_a_2_5 /= "111001010111110100100010011" OR uut_a_3_0 /= "111111110101010110101110000" OR uut_a_3_1 /= "000000111010100011000011000" OR uut_a_3_2 /= "001000011001100100101101000" OR uut_a_3_3 /= "000000000011100111001000000" OR uut_a_3_4 /= "111111101100001000110100000" OR uut_a_3_5 /= "111101001001101000001100000" OR uut_a_4_0 /= "000000000000111010100011000" OR uut_a_4_1 /= "111111111010111101111111001" OR uut_a_4_2 /= "111111010001110011010110001" OR uut_a_4_3 /= "111111111111101100001000110" OR uut_a_4_4 /= "000000000001101101001111100" OR uut_a_4_5 /= "000000001111101011000010111" OR uut_a_5_0 /= "000000001000011001100100101" OR uut_a_5_1 /= "111111010001110011010110001" OR uut_a_5_2 /= "111001010111110100100010011" OR uut_a_5_3 /= "111111111101001001101000001" OR uut_a_5_4 /= "000000001111101011000010111" OR uut_a_5_5 /= "000010001111111001110010100" THEN
              FAIL <= '1';
              FAIL_NUM <= "00011110";
              state <= "11111101";
            ELSE
              state <= "00101100";
            END IF;
            uut_rst <= '0';
          WHEN "00101100" =>
            uut_coord_shift <= "0111";
            uut_x <= "000010010100";
            uut_y <= "111110111101";
            uut_fx <= "1011010011";
            uut_fy <= "1001011001";
            uut_ft <= "0100010110";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000011010011001010000100" OR uut_a_0_1 /= "101000111001111001100100000" OR uut_a_0_2 /= "110101011110111011111011010" OR uut_a_0_3 /= "111111111111101010001101000" OR uut_a_0_4 /= "000000010011000100101000000" OR uut_a_0_5 /= "000000001000101011110100100" OR uut_a_1_0 /= "111111101000111001111001100" OR uut_a_1_1 /= "010100001101010101101000100" OR uut_a_1_2 /= "001001001100111011100100001" OR uut_a_1_3 /= "000000000000010011000100101" OR uut_a_1_4 /= "111111101111010011111101000" OR uut_a_1_5 /= "111111111000011001101010000" OR uut_a_2_0 /= "111111110101011110111011111" OR uut_a_2_1 /= "001001001100111011100100001" OR uut_a_2_2 /= "000100001100001011000111111" OR uut_a_2_3 /= "000000000000001000101011110" OR uut_a_2_4 /= "111111111000011001101010000" OR uut_a_2_5 /= "111111111100100010100010100" OR uut_a_3_0 /= "111111111111101010001101000" OR uut_a_3_1 /= "000000010011000100101000000" OR uut_a_3_2 /= "000000001000101011110100100" OR uut_a_3_3 /= "000000000000000000010010000" OR uut_a_3_4 /= "111111111111110000010000000" OR uut_a_3_5 /= "111111111111111000110101000" OR uut_a_4_0 /= "000000000000010011000100101" OR uut_a_4_1 /= "111111101111010011111101000" OR uut_a_4_2 /= "111111111000011001101010000" OR uut_a_4_3 /= "111111111111111111110000010" OR uut_a_4_4 /= "000000000000001101110010000" OR uut_a_4_5 /= "000000000000000110010001101" OR uut_a_5_0 /= "000000000000001000101011110" OR uut_a_5_1 /= "111111111000011001101010000" OR uut_a_5_2 /= "111111111100100010100010100" OR uut_a_5_3 /= "111111111111111111111000110" OR uut_a_5_4 /= "000000000000000110010001101" OR uut_a_5_5 /= "000000000000000010110110111" THEN
              FAIL <= '1';
              FAIL_NUM <= "00011111";
              state <= "11111101";
            ELSE
              state <= "00101101";
            END IF;
            uut_rst <= '0';
          WHEN "00101101" =>
            uut_coord_shift <= "0111";
            uut_x <= "111101101010";
            uut_y <= "111111000111";
            uut_fx <= "0000110101";
            uut_fy <= "1011101010";
            uut_ft <= "0010010001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000010110011101110100100" OR uut_a_0_1 /= "000101110010101100000010010" OR uut_a_0_2 /= "101101101111110001010110000" OR uut_a_0_3 /= "111111110001001000001010000" OR uut_a_0_4 /= "111100001010100110100101000" OR uut_a_0_5 /= "001100000101010111111000000" OR uut_a_1_0 /= "000000000101110010101100000" OR uut_a_1_1 /= "000001011111100100010110100" OR uut_a_1_2 /= "111011010010110100001110001" OR uut_a_1_3 /= "111111111100001010100110100" OR uut_a_1_4 /= "111111000000101110111100100" OR uut_a_1_5 /= "000011000111011000101001111" OR uut_a_2_0 /= "111111101101101111110001010" OR uut_a_2_1 /= "111011010010110100001110001" OR uut_a_2_2 /= "001110110101001011111010001" OR uut_a_2_3 /= "000000001100000101010111111" OR uut_a_2_4 /= "000011000111011000101001111" OR uut_a_2_5 /= "110110001011101000100110100" OR uut_a_3_0 /= "111111110001001000001010000" OR uut_a_3_1 /= "111100001010100110100101000" OR uut_a_3_2 /= "001100000101010111111000000" OR uut_a_3_3 /= "000000001001110110001000000" OR uut_a_3_4 /= "000010100010011101000100000" OR uut_a_3_5 /= "111000000000000001100000000" OR uut_a_4_0 /= "111111111100001010100110100" OR uut_a_4_1 /= "111111000000101110111100100" OR uut_a_4_2 /= "000011000111011000101001111" OR uut_a_4_3 /= "000000000010100010011101000" OR uut_a_4_4 /= "000000101001111000011111100" OR uut_a_4_5 /= "111101111100000000011000110" OR uut_a_5_0 /= "000000001100000101010111111" OR uut_a_5_1 /= "000011000111011000101001111" OR uut_a_5_2 /= "110110001011101000100110100" OR uut_a_5_3 /= "111111111000000000000001100" OR uut_a_5_4 /= "111101111100000000011000110" OR uut_a_5_5 /= "000110011111111110110010000" THEN
              FAIL <= '1';
              FAIL_NUM <= "00100000";
              state <= "11111101";
            ELSE
              state <= "00101110";
            END IF;
            uut_rst <= '0';
          WHEN "00101110" =>
            uut_coord_shift <= "0111";
            uut_x <= "111111111001";
            uut_y <= "111101001110";
            uut_fx <= "0100100001";
            uut_fy <= "1001100111";
            uut_ft <= "1100101101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000001101100111100010000" OR uut_a_0_1 /= "000000110110011110001000000" OR uut_a_0_2 /= "110101010111000111011100000" OR uut_a_0_3 /= "111111111001001110110110000" OR uut_a_0_4 /= "111111100100111011011000000" OR uut_a_0_5 /= "000101010010011001110100000" OR uut_a_1_0 /= "000000000000110110011110001" OR uut_a_1_1 /= "000000000011011001111000100" OR uut_a_1_2 /= "111111010101011100011101110" OR uut_a_1_3 /= "111111111111100100111011011" OR uut_a_1_4 /= "111111111110010011101101100" OR uut_a_1_5 /= "000000010101001001100111010" OR uut_a_2_0 /= "111111110101010111000111011" OR uut_a_2_1 /= "111111010101011100011101110" OR uut_a_2_2 /= "001000010011111100001100001" OR uut_a_2_3 /= "000000000101010010011001110" OR uut_a_2_4 /= "000000010101001001100111010" OR uut_a_2_5 /= "111011110111100111110101011" OR uut_a_3_0 /= "111111111001001110110110000" OR uut_a_3_1 /= "111111100100111011011000000" OR uut_a_3_2 /= "000101010010011001110100000" OR uut_a_3_3 /= "000000000011010111010010000" OR uut_a_3_4 /= "000000001101011101001000000" OR uut_a_3_5 /= "111101010111110011111100000" OR uut_a_4_0 /= "111111111111100100111011011" OR uut_a_4_1 /= "111111111110010011101101100" OR uut_a_4_2 /= "000000010101001001100111010" OR uut_a_4_3 /= "000000000000001101011101001" OR uut_a_4_4 /= "000000000000110101110100100" OR uut_a_4_5 /= "111111110101011111001111110" OR uut_a_5_0 /= "000000000101010010011001110" OR uut_a_5_1 /= "000000010101001001100111010" OR uut_a_5_2 /= "111011110111100111110101011" OR uut_a_5_3 /= "111111111101010111110011111" OR uut_a_5_4 /= "111111110101011111001111110" OR uut_a_5_5 /= "000010000011011001011011001" THEN
              FAIL <= '1';
              FAIL_NUM <= "00100001";
              state <= "11111101";
            ELSE
              state <= "00101111";
            END IF;
            uut_rst <= '0';
          WHEN "00101111" =>
            uut_coord_shift <= "0111";
            uut_x <= "111101111010";
            uut_y <= "000000001111";
            uut_fx <= "1001011110";
            uut_fy <= "1110011111";
            uut_ft <= "1001101011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000011010000011100010000" OR uut_a_0_1 /= "001100110100101111001111000" OR uut_a_0_2 /= "100110100011100011010011000" OR uut_a_0_3 /= "111111110110010011001100000" OR uut_a_0_4 /= "111011001110011100011010000" OR uut_a_0_5 /= "001001011110010000110010000" OR uut_a_1_0 /= "000000001100110100101111001" OR uut_a_1_1 /= "000110010011111101001111111" OR uut_a_1_2 /= "110011011110011111110111110" OR uut_a_1_3 /= "111111111011001110011100011" OR uut_a_1_4 /= "111101101001100110111110110" OR uut_a_1_5 /= "000100101010011001010000100" OR uut_a_2_0 /= "111111100110100011100011010" OR uut_a_2_1 /= "110011011110011111110111110" OR uut_a_2_2 /= "011000110110010010000001111" OR uut_a_2_3 /= "000000001001011110010000110" OR uut_a_2_4 /= "000100101010011001010000100" OR uut_a_2_5 /= "110110101111111100100111001" OR uut_a_3_0 /= "111111110110010011001100000" OR uut_a_3_1 /= "111011001110011100011010000" OR uut_a_3_2 /= "001001011110010000110010000" OR uut_a_3_3 /= "000000000011100111001000000" OR uut_a_3_4 /= "000001110001110000011100000" OR uut_a_3_5 /= "111100011110010010101100000" OR uut_a_4_0 /= "111111111011001110011100011" OR uut_a_4_1 /= "111101101001100110111110110" OR uut_a_4_2 /= "000100101010011001010000100" OR uut_a_4_3 /= "000000000001110001110000011" OR uut_a_4_4 /= "000000110111111111010101110" OR uut_a_4_5 /= "111110010000111010001100101" OR uut_a_5_0 /= "000000001001011110010000110" OR uut_a_5_1 /= "000100101010011001010000100" OR uut_a_5_2 /= "110110101111111100100111001" OR uut_a_5_3 /= "111111111100011110010010101" OR uut_a_5_4 /= "111110010000111010001100101" OR uut_a_5_5 /= "000011011100011010110000000" THEN
              FAIL <= '1';
              FAIL_NUM <= "00100010";
              state <= "11111101";
            ELSE
              state <= "00110000";
            END IF;
            uut_rst <= '0';
          WHEN "00110000" =>
            uut_coord_shift <= "0111";
            uut_x <= "111100111010";
            uut_y <= "000010010001";
            uut_fx <= "1100101011";
            uut_fy <= "0001101010";
            uut_ft <= "0111011100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000101011111001000000" OR uut_a_0_1 /= "000000010000011101011000000" OR uut_a_0_2 /= "000010011111000110101000000" OR uut_a_0_3 /= "000000000111011101000000000" OR uut_a_0_4 /= "000000010110010111000000000" OR uut_a_0_5 /= "000011011000001001000000000" OR uut_a_1_0 /= "000000000000010000011101011" OR uut_a_1_1 /= "000000000000110001011000001" OR uut_a_1_2 /= "000000000111011101010011111" OR uut_a_1_3 /= "000000000000010110010111000" OR uut_a_1_4 /= "000000000001000011000101000" OR uut_a_1_5 /= "000000001010001000011011000" OR uut_a_2_0 /= "000000000010011111000110101" OR uut_a_2_1 /= "000000000111011101010011111" OR uut_a_2_2 /= "000001001000000110000000001" OR uut_a_2_3 /= "000000000011011000001001000" OR uut_a_2_4 /= "000000001010001000011011000" OR uut_a_2_5 /= "000001100001111100000101000" OR uut_a_3_0 /= "000000000111011101000000000" OR uut_a_3_1 /= "000000010110010111000000000" OR uut_a_3_2 /= "000011011000001001000000000" OR uut_a_3_3 /= "000000001010001000000000000" OR uut_a_3_4 /= "000000011110011000000000000" OR uut_a_3_5 /= "000100100101101000000000000" OR uut_a_4_0 /= "000000000000010110010111000" OR uut_a_4_1 /= "000000000001000011000101000" OR uut_a_4_2 /= "000000001010001000011011000" OR uut_a_4_3 /= "000000000000011110011000000" OR uut_a_4_4 /= "000000000001011011001000000" OR uut_a_4_5 /= "000000001101110000111000000" OR uut_a_5_0 /= "000000000011011000001001000" OR uut_a_5_1 /= "000000001010001000011011000" OR uut_a_5_2 /= "000001100001111100000101000" OR uut_a_5_3 /= "000000000100100101101000000" OR uut_a_5_4 /= "000000001101110000111000000" OR uut_a_5_5 /= "000010000101000011001000000" THEN
              FAIL <= '1';
              FAIL_NUM <= "00100011";
              state <= "11111101";
            ELSE
              state <= "00110001";
            END IF;
            uut_rst <= '0';
          WHEN "00110001" =>
            uut_coord_shift <= "0111";
            uut_x <= "111111011110";
            uut_y <= "000001100011";
            uut_fx <= "0100001000";
            uut_fy <= "1110111011";
            uut_ft <= "0010011111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001010111110010000" OR uut_a_0_1 /= "000000100001100110101001000" OR uut_a_0_2 /= "000000001001100110011110000" OR uut_a_0_3 /= "000000000101110011110101000" OR uut_a_0_4 /= "000010001110010101110010100" OR uut_a_0_5 /= "000000101000101010110011000" OR uut_a_1_0 /= "000000000000100001100110101" OR uut_a_1_1 /= "000000001100110111010010101" OR uut_a_1_2 /= "000000000011101011001110011" OR uut_a_1_3 /= "000000000010001110010101110" OR uut_a_1_4 /= "000000110110011111010101110" OR uut_a_1_5 /= "000000001111100100011000100" OR uut_a_2_0 /= "000000000000001001100110011" OR uut_a_2_1 /= "000000000011101011001110011" OR uut_a_2_2 /= "000000000001000011001101010" OR uut_a_2_3 /= "000000000000101000101010110" OR uut_a_2_4 /= "000000001111100100011000100" OR uut_a_2_5 /= "000000000100011100101011100" OR uut_a_3_0 /= "000000000101110011110101000" OR uut_a_3_1 /= "000010001110010101110010100" OR uut_a_3_2 /= "000000101000101010110011000" OR uut_a_3_3 /= "000000011000100111000000100" OR uut_a_3_4 /= "001001011010111011101100010" OR uut_a_3_5 /= "000010101100010001000011100" OR uut_a_4_0 /= "000000000010001110010101110" OR uut_a_4_1 /= "000000110110011111010101110" OR uut_a_4_2 /= "000000001111100100011000100" OR uut_a_4_3 /= "000000001001011010111011101" OR uut_a_4_4 /= "000011100110110011110110011" OR uut_a_4_5 /= "000001000001111100100001110" OR uut_a_5_0 /= "000000000000101000101010110" OR uut_a_5_1 /= "000000001111100100011000100" OR uut_a_5_2 /= "000000000100011100101011100" OR uut_a_5_3 /= "000000000010101100010001000" OR uut_a_5_4 /= "000001000001111100100001110" OR uut_a_5_5 /= "000000010010110101110111011" THEN
              FAIL <= '1';
              FAIL_NUM <= "00100100";
              state <= "11111101";
            ELSE
              state <= "00110010";
            END IF;
            uut_rst <= '0';
          WHEN "00110010" =>
            uut_coord_shift <= "0111";
            uut_x <= "111100111001";
            uut_y <= "000011011110";
            uut_fx <= "1011000000";
            uut_fy <= "1100010001";
            uut_ft <= "0100110001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000111011100101000100" OR uut_a_0_1 /= "111101100111010101000001110" OR uut_a_0_2 /= "000001100100100010100010110" OR uut_a_0_3 /= "111111110011110010011110100" OR uut_a_0_4 /= "000011111010010101001110110" OR uut_a_0_5 /= "111101011011001001011011110" OR uut_a_1_0 /= "111111111101100111010101000" OR uut_a_1_1 /= "000000110000111001110000111" OR uut_a_1_2 /= "111111011111110010111011110" OR uut_a_1_3 /= "000000000011111010010101001" OR uut_a_1_4 /= "111110101111110100001100110" OR uut_a_1_5 /= "000000110100110011011110100" OR uut_a_2_0 /= "000000000001100100100010100" OR uut_a_2_1 /= "111111011111110010111011110" OR uut_a_2_2 /= "000000010101001101010010010" OR uut_a_2_3 /= "111111111101011011001001011" OR uut_a_2_4 /= "000000110100110011011110100" OR uut_a_2_5 /= "111111011101001110011111010" OR uut_a_3_0 /= "111111110011110010011110100" OR uut_a_3_1 /= "000011111010010101001110110" OR uut_a_3_2 /= "111101011011001001011011110" OR uut_a_3_3 /= "000000010100000001011100100" OR uut_a_3_4 /= "111001100101100010010111110" OR uut_a_3_5 /= "000100001110010011100000110" OR uut_a_4_0 /= "000000000011111010010101001" OR uut_a_4_1 /= "111110101111110100001100110" OR uut_a_4_2 /= "000000110100110011011110100" OR uut_a_4_3 /= "111111111001100101100010010" OR uut_a_4_4 /= "000010000011011110011111011" OR uut_a_4_5 /= "111110101001011010110000000" OR uut_a_5_0 /= "111111111101011011001001011" OR uut_a_5_1 /= "000000110100110011011110100" OR uut_a_5_2 /= "111111011101001110011111010" OR uut_a_5_3 /= "000000000100001110010011100" OR uut_a_5_4 /= "111110101001011010110000000" OR uut_a_5_5 /= "000000111001000001000111011" THEN
              FAIL <= '1';
              FAIL_NUM <= "00100101";
              state <= "11111101";
            ELSE
              state <= "00110011";
            END IF;
            uut_rst <= '0';
          WHEN "00110011" =>
            uut_coord_shift <= "0111";
            uut_x <= "111111111010";
            uut_y <= "000010001001";
            uut_fx <= "1110010110";
            uut_fy <= "1100010111";
            uut_ft <= "1000100110";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000010011100010000000000" OR uut_a_0_1 /= "000001110101001100000000000" OR uut_a_0_2 /= "111111100010101101000000000" OR uut_a_0_3 /= "000000001110111100010000000" OR uut_a_0_4 /= "000001011001101001100000000" OR uut_a_0_5 /= "111111101001100101101000000" OR uut_a_1_0 /= "000000000001110101001100000" OR uut_a_1_1 /= "000000001010111111001000000" OR uut_a_1_2 /= "111111111101010000001110000" OR uut_a_1_3 /= "000000000001011001101001100" OR uut_a_1_4 /= "000000001000011001111001000" OR uut_a_1_5 /= "111111111101111001100001110" OR uut_a_2_0 /= "111111111111100010101101000" OR uut_a_2_1 /= "111111111101010000001110000" OR uut_a_2_2 /= "000000000000101011111100100" OR uut_a_2_3 /= "111111111111101001100101101" OR uut_a_2_4 /= "111111111101111001100001110" OR uut_a_2_5 /= "000000000000100001100111100" OR uut_a_3_0 /= "000000001110111100010000000" OR uut_a_3_1 /= "000001011001101001100000000" OR uut_a_3_2 /= "111111101001100101101000000" OR uut_a_3_3 /= "000000001011011011100010000" OR uut_a_3_4 /= "000001000100100101001100000" OR uut_a_3_5 /= "111111101110110110101101000" OR uut_a_4_0 /= "000000000001011001101001100" OR uut_a_4_1 /= "000000001000011001111001000" OR uut_a_4_2 /= "111111111101111001100001110" OR uut_a_4_3 /= "000000000001000100100101001" OR uut_a_4_4 /= "000000000110011011011111001" OR uut_a_4_5 /= "111111111110011001001000001" OR uut_a_5_0 /= "111111111111101001100101101" OR uut_a_5_1 /= "111111111101111001100001110" OR uut_a_5_2 /= "000000000000100001100111100" OR uut_a_5_3 /= "111111111111101110110110101" OR uut_a_5_4 /= "111111111110011001001000001" OR uut_a_5_5 /= "000000000000011001101101111" THEN
              FAIL <= '1';
              FAIL_NUM <= "00100110";
              state <= "11111101";
            ELSE
              state <= "00110100";
            END IF;
            uut_rst <= '0';
          WHEN "00110100" =>
            uut_coord_shift <= "0111";
            uut_x <= "000001011000";
            uut_y <= "111111011100";
            uut_fx <= "1111001111";
            uut_fy <= "0001110000";
            uut_ft <= "1000111101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000010101101000101100100" OR uut_a_0_1 /= "101100101110110000010111100" OR uut_a_0_2 /= "101101100100110110000110110" OR uut_a_0_3 /= "111111110000010001100011000" OR uut_a_0_4 /= "001110000000010111110101000" OR uut_a_0_5 /= "001101011001000011101100100" OR uut_a_1_0 /= "111111101100101110110000010" OR uut_a_1_1 /= "010001001010010110111011000" OR uut_a_1_2 /= "010000011010001011110011111" OR uut_a_1_3 /= "000000001110000000010111110" OR uut_a_1_4 /= "110011100001101010110001110" OR uut_a_1_5 /= "110100000100101011101101010" OR uut_a_2_0 /= "111111101101100100110110000" OR uut_a_2_1 /= "010000011010001011110011111" OR uut_a_2_2 /= "001111101100000111111011010" OR uut_a_2_3 /= "000000001101011001000011101" OR uut_a_2_4 /= "110100000100101011101101010" OR uut_a_2_5 /= "110100100110001010010110100" OR uut_a_3_0 /= "111111110000010001100011000" OR uut_a_3_1 /= "001110000000010111110101000" OR uut_a_3_2 /= "001101011001000011101100100" OR uut_a_3_3 /= "000000001011011011100010000" OR uut_a_3_4 /= "110101110100011110101110000" OR uut_a_3_5 /= "110110010001000011100011000" OR uut_a_4_0 /= "000000001110000000010111110" OR uut_a_4_1 /= "110011100001101010110001110" OR uut_a_4_2 /= "110100000100101011101101010" OR uut_a_4_3 /= "111111110101110100011110101" OR uut_a_4_4 /= "001001000100010000101001000" OR uut_a_4_5 /= "001000101010110011110101110" OR uut_a_5_0 /= "000000001101011001000011101" OR uut_a_5_1 /= "110100000100101011101101010" OR uut_a_5_2 /= "110100100110001010010110100" OR uut_a_5_3 /= "111111110110010001000011100" OR uut_a_5_4 /= "001000101010110011110101110" OR uut_a_5_5 /= "001000010010011110011110101" THEN
              FAIL <= '1';
              FAIL_NUM <= "00100111";
              state <= "11111101";
            ELSE
              state <= "00110101";
            END IF;
            uut_rst <= '0';
          WHEN "00110101" =>
            uut_coord_shift <= "0111";
            uut_x <= "111110100010";
            uut_y <= "000010001011";
            uut_fx <= "0011001001";
            uut_fy <= "1010000000";
            uut_ft <= "1010000101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000011001011000100000" OR uut_a_0_1 /= "000010010101000111111100000" OR uut_a_0_2 /= "111011010101110000001000000" OR uut_a_0_3 /= "111111111010011100101001000" OR uut_a_0_4 /= "111011111011000010000111000" OR uut_a_0_5 /= "001000001001111011110010000" OR uut_a_1_0 /= "000000000001001010100011111" OR uut_a_1_1 /= "000000110110110000011010100" OR uut_a_1_2 /= "111110010010011111001010111" OR uut_a_1_3 /= "111111111101111101100001000" OR uut_a_1_4 /= "111110100000001011010001100" OR uut_a_1_5 /= "000010111111101001011100110" OR uut_a_2_0 /= "111111111101101010111000000" OR uut_a_2_1 /= "111110010010011111001010111" OR uut_a_2_2 /= "000011011011000001101010001" OR uut_a_2_3 /= "000000000100000100111101111" OR uut_a_2_4 /= "000010111111101001011100110" OR uut_a_2_5 /= "111010000000101101000110010" OR uut_a_3_0 /= "111111111010011100101001000" OR uut_a_3_1 /= "111011111011000010000111000" OR uut_a_3_2 /= "001000001001111011110010000" OR uut_a_3_3 /= "000000001001101101111000010" OR uut_a_3_4 /= "000111001000101100010011110" OR uut_a_3_5 /= "110001101110100111011000100" OR uut_a_4_0 /= "111111111101111101100001000" OR uut_a_4_1 /= "111110100000001011010001100" OR uut_a_4_2 /= "000010111111101001011100110" OR uut_a_4_3 /= "000000000011100100010110001" OR uut_a_4_4 /= "000010100111101100010001010" OR uut_a_4_5 /= "111010110000100111011101011" OR uut_a_5_0 /= "000000000100000100111101111" OR uut_a_5_1 /= "000010111111101001011100110" OR uut_a_5_2 /= "111010000000101101000110010" OR uut_a_5_3 /= "111111111000110111010011101" OR uut_a_5_4 /= "111010110000100111011101011" OR uut_a_5_5 /= "001010011110110001000101000" THEN
              FAIL <= '1';
              FAIL_NUM <= "00101000";
              state <= "11111101";
            ELSE
              state <= "00110110";
            END IF;
            uut_rst <= '0';
          WHEN "00110110" =>
            uut_coord_shift <= "0111";
            uut_x <= "111100110000";
            uut_y <= "111100000101";
            uut_fx <= "1110110001";
            uut_fy <= "0010011111";
            uut_ft <= "0011100100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001100001100001000" OR uut_a_0_1 /= "000000110110110110100100000" OR uut_a_0_2 /= "111110111101101110000100100" OR uut_a_0_3 /= "000000000010011101011000100" OR uut_a_0_4 /= "000001011000100001110010000" OR uut_a_0_5 /= "111110010101000001110110010" OR uut_a_1_0 /= "000000000000011011011011010" OR uut_a_1_1 /= "000000001111011011010110001" OR uut_a_1_2 /= "111111101101010110111101010" OR uut_a_1_3 /= "000000000000101100010000111" OR uut_a_1_4 /= "000000011000111001100000000" OR uut_a_1_5 /= "111111100001111010100001010" OR uut_a_2_0 /= "111111111111011110110111000" OR uut_a_2_1 /= "111111101101010110111101010" OR uut_a_2_2 /= "000000010110100001100101111" OR uut_a_2_3 /= "111111111111001010100000111" OR uut_a_2_4 /= "111111100001111010100001010" OR uut_a_2_5 /= "000000100100010110100111110" OR uut_a_3_0 /= "000000000010011101011000100" OR uut_a_3_1 /= "000001011000100001110010000" OR uut_a_3_2 /= "111110010101000001110110010" OR uut_a_3_3 /= "000000000011111110000000010" OR uut_a_3_4 /= "000010001110111000001001000" OR uut_a_3_5 /= "111101010011010110110101001" OR uut_a_4_0 /= "000000000000101100010000111" OR uut_a_4_1 /= "000000011000111001100000000" OR uut_a_4_2 /= "111111100001111010100001010" OR uut_a_4_3 /= "000000000001000111011100000" OR uut_a_4_4 /= "000000101000001011110010100" OR uut_a_4_5 /= "111111001111011100011010111" OR uut_a_5_0 /= "111111111111001010100000111" OR uut_a_5_1 /= "111111100001111010100001010" OR uut_a_5_2 /= "000000100100010110100111110" OR uut_a_5_3 /= "111111111110101001101011011" OR uut_a_5_4 /= "111111001111011100011010111" OR uut_a_5_5 /= "000000111010101010111111011" THEN
              FAIL <= '1';
              FAIL_NUM <= "00101001";
              state <= "11111101";
            ELSE
              state <= "00110111";
            END IF;
            uut_rst <= '0';
          WHEN "00110111" =>
            uut_coord_shift <= "0111";
            uut_x <= "000000001111";
            uut_y <= "111100111000";
            uut_fx <= "0010000111";
            uut_fy <= "1010000010";
            uut_ft <= "1010001010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000011100010111000010" OR uut_a_0_1 /= "000011011000001111100111010" OR uut_a_0_2 /= "111100010000101101101011001" OR uut_a_0_3 /= "000000000111000101110000100" OR uut_a_0_4 /= "000110110000011111001110100" OR uut_a_0_5 /= "111000100001011011010110010" OR uut_a_1_0 /= "000000000001101100000111110" OR uut_a_1_1 /= "000001100111000011011100001" OR uut_a_1_2 /= "111110001101111101110001000" OR uut_a_1_3 /= "000000000011011000001111100" OR uut_a_1_4 /= "000011001110000110111000011" OR uut_a_1_5 /= "111100011011111011100010000" OR uut_a_2_0 /= "111111111110001000010110110" OR uut_a_2_1 /= "111110001101111101110001000" OR uut_a_2_2 /= "000001111110001011111010100" OR uut_a_2_3 /= "111111111100010000101101101" OR uut_a_2_4 /= "111100011011111011100010000" OR uut_a_2_5 /= "000011111100010111110101000" OR uut_a_3_0 /= "000000000111000101110000100" OR uut_a_3_1 /= "000110110000011111001110100" OR uut_a_3_2 /= "111000100001011011010110010" OR uut_a_3_3 /= "000000001110001011100001000" OR uut_a_3_4 /= "001101100000111110011101000" OR uut_a_3_5 /= "110001000010110110101100100" OR uut_a_4_0 /= "000000000011011000001111100" OR uut_a_4_1 /= "000011001110000110111000011" OR uut_a_4_2 /= "111100011011111011100010000" OR uut_a_4_3 /= "000000000110110000011111001" OR uut_a_4_4 /= "000110011100001101110000110" OR uut_a_4_5 /= "111000110111110111000100001" OR uut_a_5_0 /= "111111111100010000101101101" OR uut_a_5_1 /= "111100011011111011100010000" OR uut_a_5_2 /= "000011111100010111110101000" OR uut_a_5_3 /= "111111111000100001011011010" OR uut_a_5_4 /= "111000110111110111000100001" OR uut_a_5_5 /= "000111111000101111101010000" THEN
              FAIL <= '1';
              FAIL_NUM <= "00101010";
              state <= "11111101";
            ELSE
              state <= "00111000";
            END IF;
            uut_rst <= '0';
          WHEN "00111000" =>
            uut_coord_shift <= "0111";
            uut_x <= "111100110011";
            uut_y <= "111101001001";
            uut_fx <= "1010101100";
            uut_fy <= "1011001001";
            uut_ft <= "1101000101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001000110001001000" OR uut_a_0_1 /= "111110001100011000001010100" OR uut_a_0_2 /= "111111011010101111001110000" OR uut_a_0_3 /= "111111111110011101000100100" OR uut_a_0_4 /= "000010100011000101000101010" OR uut_a_0_5 /= "000000110100100011100111000" OR uut_a_1_0 /= "111111111111000110001100000" OR uut_a_1_1 /= "000001011111010011000101010" OR uut_a_1_2 /= "000000011110101101100101001" OR uut_a_1_3 /= "000000000001010001100010100" OR uut_a_1_4 /= "111101111001100101100011111" OR uut_a_1_5 /= "111111010100101011101001100" OR uut_a_2_0 /= "111111111111101101010111100" OR uut_a_2_1 /= "000000011110101101100101001" OR uut_a_2_2 /= "000000001001111001011101010" OR uut_a_2_3 /= "000000000000011010010001110" OR uut_a_2_4 /= "111111010100101011101001100" OR uut_a_2_5 /= "111111110010000010100010101" OR uut_a_3_0 /= "111111111110011101000100100" OR uut_a_3_1 /= "000010100011000101000101010" OR uut_a_3_2 /= "000000110100100011100111000" OR uut_a_3_3 /= "000000000010001011100010010" OR uut_a_3_4 /= "111100011001111111000010101" OR uut_a_3_5 /= "111110110101110111110011100" OR uut_a_4_0 /= "000000000001010001100010100" OR uut_a_4_1 /= "111101111001100101100011111" OR uut_a_4_2 /= "111111010100101011101001100" OR uut_a_4_3 /= "111111111110001100111111100" OR uut_a_4_4 /= "000010111101100101010010100" OR uut_a_4_5 /= "000000111101000110010000010" OR uut_a_5_0 /= "000000000000011010010001110" OR uut_a_5_1 /= "111111010100101011101001100" OR uut_a_5_2 /= "111111110010000010100010101" OR uut_a_5_3 /= "111111111111011010111011111" OR uut_a_5_4 /= "000000111101000110010000010" OR uut_a_5_5 /= "000000010011101100001011010" THEN
              FAIL <= '1';
              FAIL_NUM <= "00101011";
              state <= "11111101";
            ELSE
              state <= "00111001";
            END IF;
            uut_rst <= '0';
          WHEN "00111001" =>
            uut_coord_shift <= "0111";
            uut_x <= "111110100011";
            uut_y <= "111101110000";
            uut_fx <= "1100000001";
            uut_fy <= "0110010010";
            uut_ft <= "0011010000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000101100001111010010" OR uut_a_0_1 /= "000110011001001101010110100" OR uut_a_0_2 /= "111101000110110000000000101" OR uut_a_0_3 /= "000000000111110001010110110" OR uut_a_0_4 /= "001000111111000100010011100" OR uut_a_0_5 /= "111011111011101010100101111" OR uut_a_1_0 /= "000000000011001100100110101" OR uut_a_1_1 /= "000011101100100100101110000" OR uut_a_1_2 /= "111110010100111001110000010" OR uut_a_1_3 /= "000000000100011111100010001" OR uut_a_1_4 /= "000101001100011101011111010" OR uut_a_1_5 /= "111101101001011111100111111" OR uut_a_2_0 /= "111111111110100011011000000" OR uut_a_2_1 /= "111110010100111001110000010" OR uut_a_2_2 /= "000000110000011110111011110" OR uut_a_2_3 /= "111111111101111101110101010" OR uut_a_2_4 /= "111101101001011111100111111" OR uut_a_2_5 /= "000001000100001000100110100" OR uut_a_3_0 /= "000000000111110001010110110" OR uut_a_3_1 /= "001000111111000100010011100" OR uut_a_3_2 /= "111011111011101010100101111" OR uut_a_3_3 /= "000000001010111010111100010" OR uut_a_3_4 /= "001100101000001001101010100" OR uut_a_3_5 /= "111010010010001001011101101" OR uut_a_4_0 /= "000000000100011111100010001" OR uut_a_4_1 /= "000101001100011101011111010" OR uut_a_4_2 /= "111101101001011111100111111" OR uut_a_4_3 /= "000000000110010100000100110" OR uut_a_4_4 /= "000111010011001101100101100" OR uut_a_4_5 /= "111100101100011111011110001" OR uut_a_5_0 /= "111111111101111101110101010" OR uut_a_5_1 /= "111101101001011111100111111" OR uut_a_5_2 /= "000001000100001000100110100" OR uut_a_5_3 /= "111111111101001001000100101" OR uut_a_5_4 /= "111100101100011111011110001" OR uut_a_5_5 /= "000001011111110000000001011" THEN
              FAIL <= '1';
              FAIL_NUM <= "00101100";
              state <= "11111101";
            ELSE
              state <= "00111010";
            END IF;
            uut_rst <= '0';
          WHEN "00111010" =>
            uut_coord_shift <= "0111";
            uut_x <= "000000011100";
            uut_y <= "111101011111";
            uut_fx <= "1011011001";
            uut_fy <= "1001001111";
            uut_ft <= "0110101000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000001010111110010" OR uut_a_0_1 /= "111111110011001001000011010" OR uut_a_0_2 /= "111111111011000111010001111" OR uut_a_0_3 /= "111111111111000110011100100" OR uut_a_0_4 /= "000001000011011100100110100" OR uut_a_0_5 /= "000000011001101000010011110" OR uut_a_1_0 /= "111111111111111001100100100" OR uut_a_1_1 /= "000000000111100010001100100" OR uut_a_1_2 /= "000000000010110111001111000" OR uut_a_1_3 /= "000000000000100001101110010" OR uut_a_1_4 /= "111111011000011110101111011" OR uut_a_1_5 /= "111111110000111110111000011" OR uut_a_2_0 /= "111111111111111101100011101" OR uut_a_2_1 /= "000000000010110111001111000" OR uut_a_2_2 /= "000000000001000101101000010" OR uut_a_2_3 /= "000000000000001100110100001" OR uut_a_2_4 /= "111111110000111110111000011" OR uut_a_2_5 /= "111111111010010010110001100" OR uut_a_3_0 /= "111111111111000110011100100" OR uut_a_3_1 /= "000001000011011100100110100" OR uut_a_3_2 /= "000000011001101000010011110" OR uut_a_3_3 /= "000000000100101101111001000" OR uut_a_3_4 /= "111010011110001110001101000" OR uut_a_3_5 /= "111101111001100100000111100" OR uut_a_4_0 /= "000000000000100001101110010" OR uut_a_4_1 /= "111111011000011110101111011" OR uut_a_4_2 /= "111111110000111110111000011" OR uut_a_4_3 /= "111111111101001111000111000" OR uut_a_4_4 /= "000011001111010010101011011" OR uut_a_4_5 /= "000001001110110001010101100" OR uut_a_5_0 /= "000000000000001100110100001" OR uut_a_5_1 /= "111111110000111110111000011" OR uut_a_5_2 /= "111111111010010010110001100" OR uut_a_5_3 /= "111111111110111100110010000" OR uut_a_5_4 /= "000001001110110001010101100" OR uut_a_5_5 /= "000000011101111011101101010" THEN
              FAIL <= '1';
              FAIL_NUM <= "00101101";
              state <= "11111101";
            ELSE
              state <= "00111011";
            END IF;
            uut_rst <= '0';
          WHEN "00111011" =>
            uut_coord_shift <= "0111";
            uut_x <= "000001101001";
            uut_y <= "000000011101";
            uut_fx <= "1101000001";
            uut_fy <= "1010101010";
            uut_ft <= "0001111101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000101000110010000010" OR uut_a_0_1 /= "111111101110001010000111001" OR uut_a_0_2 /= "111000111010010011011001110" OR uut_a_0_3 /= "111111111000110010010001110" OR uut_a_0_4 /= "000000011001010000000001111" OR uut_a_0_5 /= "001010000010000101010100010" OR uut_a_1_0 /= "111111111111110111000101000" OR uut_a_1_1 /= "000000000000011111001110010" OR uut_a_1_2 /= "000000001100011001111110000" OR uut_a_1_3 /= "000000000000001100101000000" OR uut_a_1_4 /= "111111111111010011110011111" OR uut_a_1_5 /= "111111101110011100010110101" OR uut_a_2_0 /= "111111111100011101001001101" OR uut_a_2_1 /= "000000001100011001111110000" OR uut_a_2_2 /= "000100111011011101100000100" OR uut_a_2_3 /= "000000000101000001000010101" OR uut_a_2_4 /= "111111101110011100010110101" OR uut_a_2_5 /= "111001000001100011010011011" OR uut_a_3_0 /= "111111111000110010010001110" OR uut_a_3_1 /= "000000011001010000000001111" OR uut_a_3_2 /= "001010000010000101010100010" OR uut_a_3_3 /= "000000001010001101011100010" OR uut_a_3_4 /= "111111011100010000111101001" OR uut_a_3_5 /= "110001110011010011101101110" OR uut_a_4_0 /= "000000000000001100101000000" OR uut_a_4_1 /= "111111111111010011110011111" OR uut_a_4_2 /= "111111101110011100010110101" OR uut_a_4_3 /= "111111111111101110001000011" OR uut_a_4_4 /= "000000000000111110100010010" OR uut_a_4_5 /= "000000011000110110001101011" OR uut_a_5_0 /= "000000000101000001000010101" OR uut_a_5_1 /= "111111101110011100010110101" OR uut_a_5_2 /= "111001000001100011010011011" OR uut_a_5_3 /= "111111111000111001101001110" OR uut_a_5_4 /= "000000011000110110001101011" OR uut_a_5_5 /= "001001110111110100110010101" THEN
              FAIL <= '1';
              FAIL_NUM <= "00101110";
              state <= "11111101";
            ELSE
              state <= "00111100";
            END IF;
            uut_rst <= '0';
          WHEN "00111100" =>
            uut_coord_shift <= "1000";
            uut_x <= "000111110011";
            uut_y <= "111010101111";
            uut_fx <= "1100001000";
            uut_fy <= "1110010110";
            uut_ft <= "1001001100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000001010101010100001000" OR uut_a_0_1 /= "110100110101011111011101000" OR uut_a_0_2 /= "000001001111111110110111100" OR uut_a_0_3 /= "000000000010011110011000100" OR uut_a_0_4 /= "111101011010001100010110100" OR uut_a_0_5 /= "000000010010100011110111110" OR uut_a_1_0 /= "111111111010011010101111101" OR uut_a_1_1 /= "000101110110000000000010010" OR uut_a_1_2 /= "111111010110001000100101111" OR uut_a_1_3 /= "111111111110101101000110001" OR uut_a_1_4 /= "000001010110110010100010001" OR uut_a_1_5 /= "111111110110010010001110010" OR uut_a_2_0 /= "000000000000100111111111011" OR uut_a_2_1 /= "111111010110001000100101111" OR uut_a_2_2 /= "000000000100101011111011110" OR uut_a_2_3 /= "000000000000001001010001111" OR uut_a_2_4 /= "111111110110010010001110010" OR uut_a_2_5 /= "000000000001000101100110100" OR uut_a_3_0 /= "000000000010011110011000100" OR uut_a_3_1 /= "111101011010001100010110100" OR uut_a_3_2 /= "000000010010100011110111110" OR uut_a_3_3 /= "000000000000100100110000010" OR uut_a_3_4 /= "111111011001100001011111010" OR uut_a_3_5 /= "000000000100010011101001111" OR uut_a_4_0 /= "111111111110101101000110001" OR uut_a_4_1 /= "000001010110110010100010001" OR uut_a_4_2 /= "111111110110010010001110010" OR uut_a_4_3 /= "111111111111101100110000101" OR uut_a_4_4 /= "000000010100001000111110001" OR uut_a_4_5 /= "111111111101101111101101100" OR uut_a_5_0 /= "000000000000001001010001111" OR uut_a_5_1 /= "111111110110010010001110010" OR uut_a_5_2 /= "000000000001000101100110100" OR uut_a_5_3 /= "000000000000000010001001110" OR uut_a_5_4 /= "111111111101101111101101100" OR uut_a_5_5 /= "000000000000010000001001101" THEN
              FAIL <= '1';
              FAIL_NUM <= "00101111";
              state <= "11111101";
            ELSE
              state <= "00111101";
            END IF;
            uut_rst <= '0';
          WHEN "00111101" =>
            uut_coord_shift <= "1000";
            uut_x <= "000010111100";
            uut_y <= "111110011101";
            uut_fx <= "0111101110";
            uut_fy <= "1110011100";
            uut_ft <= "0001111100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000010110001001110010" OR uut_a_0_1 /= "111011101101110110111101010" OR uut_a_0_2 /= "000011001000110000101001001" OR uut_a_0_3 /= "111111111110100111110011100" OR uut_a_0_4 /= "000010001000011011010101100" OR uut_a_0_5 /= "111110011100000101110101110" OR uut_a_1_0 /= "111111111101110110111011011" OR uut_a_1_1 /= "000011010100000001111111101" OR uut_a_1_2 /= "111101100100101110011000001" OR uut_a_1_3 /= "000000000001000100001101101" OR uut_a_1_4 /= "111110010110011110110110110" OR uut_a_1_5 /= "000001001101010001011110111" OR uut_a_2_0 /= "000000000001100100011000010" OR uut_a_2_1 /= "111101100100101110011000001" OR uut_a_2_2 /= "000001110001101101100011010" OR uut_a_2_3 /= "111111111111001110000010111" OR uut_a_2_4 /= "000001001101010001011110111" OR uut_a_2_5 /= "111111000111011010010011101" OR uut_a_3_0 /= "111111111110100111110011100" OR uut_a_3_1 /= "000010001000011011010101100" OR uut_a_3_2 /= "111110011100000101110101110" OR uut_a_3_3 /= "000000000000101011111001000" OR uut_a_3_4 /= "111110111100000110110101000" OR uut_a_3_5 /= "000000110001101110000100100" OR uut_a_4_0 /= "000000000001000100001101101" OR uut_a_4_1 /= "111110010110011110110110110" OR uut_a_4_2 /= "000001001101010001011110111" OR uut_a_4_3 /= "111111111111011110000011011" OR uut_a_4_4 /= "000000110100100000101110000" OR uut_a_4_5 /= "111111011001100010110111100" OR uut_a_5_0 /= "111111111111001110000010111" OR uut_a_5_1 /= "000001001101010001011110111" OR uut_a_5_2 /= "111111000111011010010011101" OR uut_a_5_3 /= "000000000000011000110111000" OR uut_a_5_4 /= "111111011001100010110111100" OR uut_a_5_5 /= "000000011100001010010110000" THEN
              FAIL <= '1';
              FAIL_NUM <= "00110000";
              state <= "11111101";
            ELSE
              state <= "00111110";
            END IF;
            uut_rst <= '0';
          WHEN "00111110" =>
            uut_coord_shift <= "1000";
            uut_x <= "111010011111";
            uut_y <= "111110000111";
            uut_fx <= "1010100101";
            uut_fy <= "0100001000";
            uut_ft <= "0101111100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000100010000010000000" OR uut_a_0_1 /= "111110110111101011110000000" OR uut_a_0_2 /= "000011010010100100011000000" OR uut_a_0_3 /= "111111111110111000110110000" OR uut_a_0_4 /= "000000010010111001101010000" OR uut_a_0_5 /= "111111001000111101110001000" OR uut_a_1_0 /= "111111111111011011110101111" OR uut_a_1_1 /= "000000001001100110101100001" OR uut_a_1_2 /= "111111100100000010001010110" OR uut_a_1_3 /= "000000000000001001011100110" OR uut_a_1_4 /= "111111111101011111010101111" OR uut_a_1_5 /= "000000000111010011110010111" OR uut_a_2_0 /= "000000000001101001010010001" OR uut_a_2_1 /= "111111100100000010001010110" OR uut_a_2_2 /= "000001010001011011100100010" OR uut_a_2_3 /= "111111111111100100011110111" OR uut_a_2_4 /= "000000000111010011110010111" OR uut_a_2_5 /= "111111101010101101111000101" OR uut_a_3_0 /= "111111111110111000110110000" OR uut_a_3_1 /= "000000010010111001101010000" OR uut_a_3_2 /= "111111001000111101110001000" OR uut_a_3_3 /= "000000000000010010100110010" OR uut_a_3_4 /= "111111111011000011110101110" OR uut_a_3_5 /= "000000001110011000100101011" OR uut_a_4_0 /= "000000000000001001011100110" OR uut_a_4_1 /= "111111111101011111010101111" OR uut_a_4_2 /= "000000000111010011110010111" OR uut_a_4_3 /= "111111111111111101100001111" OR uut_a_4_4 /= "000000000000101001111111010" OR uut_a_4_5 /= "111111111110000101101111000" OR uut_a_5_0 /= "111111111111100100011110111" OR uut_a_5_1 /= "000000000111010011110010111" OR uut_a_5_2 /= "111111101010101101111000101" OR uut_a_5_3 /= "000000000000000111001100010" OR uut_a_5_4 /= "111111111110000101101111000" OR uut_a_5_5 /= "000000000101100100000000011" THEN
              FAIL <= '1';
              FAIL_NUM <= "00110001";
              state <= "11111101";
            ELSE
              state <= "00111111";
            END IF;
            uut_rst <= '0';
          WHEN "00111111" =>
            uut_coord_shift <= "1000";
            uut_x <= "111101101000";
            uut_y <= "000010111101";
            uut_fx <= "1100101101";
            uut_fy <= "0000011111";
            uut_ft <= "0101010100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000110010000000000000" OR uut_a_0_1 /= "110110010010001000000000000" OR uut_a_0_2 /= "001010110101110000000000000" OR uut_a_0_3 /= "000000000100101010110000000" OR uut_a_0_4 /= "111000101111100010011000000" OR uut_a_0_5 /= "001000000110001001010000000" OR uut_a_1_0 /= "111111111011001001000100000" OR uut_a_1_1 /= "000111100011011010010010000" OR uut_a_1_2 /= "110111100100101101111100000" OR uut_a_1_3 /= "111111111100010111110001001" OR uut_a_1_4 /= "000101101001000011000001110" OR uut_a_1_5 /= "111001101101001110010011110" OR uut_a_2_0 /= "000000000101011010111000000" OR uut_a_2_1 /= "110111100100101101111100000" OR uut_a_2_2 /= "001001011001100111001000000" OR uut_a_2_3 /= "000000000100000011000100101" OR uut_a_2_4 /= "111001101101001110010011110" OR uut_a_2_5 /= "000111000001010101000001011" OR uut_a_3_0 /= "000000000100101010110000000" OR uut_a_3_1 /= "111000101111100010011000000" OR uut_a_3_2 /= "001000000110001001010000000" OR uut_a_3_3 /= "000000000011011111001000010" OR uut_a_3_4 /= "111010100101000110101011001" OR uut_a_3_5 /= "000110000010111111010011110" OR uut_a_4_0 /= "111111111100010111110001001" OR uut_a_4_1 /= "000101101001000011000001110" OR uut_a_4_2 /= "111001101101001110010011110" OR uut_a_4_3 /= "111111111101010010100011010" OR uut_a_4_4 /= "000100001101101010000011111" OR uut_a_4_5 /= "111011010011001011010010011" OR uut_a_5_0 /= "000000000100000011000100101" OR uut_a_5_1 /= "111001101101001110010011110" OR uut_a_5_2 /= "000111000001010101000001011" OR uut_a_5_3 /= "000000000011000001011111101" OR uut_a_5_4 /= "111011010011001011010010011" OR uut_a_5_5 /= "000101001111100101111001101" THEN
              FAIL <= '1';
              FAIL_NUM <= "00110010";
              state <= "11111101";
            ELSE
              state <= "01000000";
            END IF;
            uut_rst <= '0';
          WHEN "01000000" =>
            uut_coord_shift <= "1000";
            uut_x <= "000001100011";
            uut_y <= "111101011000";
            uut_fx <= "1100110010";
            uut_fy <= "1111001111";
            uut_ft <= "1110110001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000101011111001000" OR uut_a_0_1 /= "111111111101111100010101000" OR uut_a_0_2 /= "000000101110111110100000100" OR uut_a_0_3 /= "000000000001100000011110100" OR uut_a_0_4 /= "111111111011011110100100100" OR uut_a_0_5 /= "000001100111010000101001010" OR uut_a_1_0 /= "111111111111111110111110001" OR uut_a_1_1 /= "000000000000000011000101100" OR uut_a_1_2 /= "111111111110111001100010001" OR uut_a_1_3 /= "111111111111111101101111010" OR uut_a_1_4 /= "000000000000000110110010001" OR uut_a_1_5 /= "111111111101100101000111000" OR uut_a_2_0 /= "000000000000010111011111010" OR uut_a_2_1 /= "111111111110111001100010001" OR uut_a_2_2 /= "000000011001001000111100111" OR uut_a_2_3 /= "000000000000110011101000010" OR uut_a_2_4 /= "111111111101100101000111000" OR uut_a_2_5 /= "000000110111010000101010000" OR uut_a_3_0 /= "000000000001100000011110100" OR uut_a_3_1 /= "111111111011011110100100100" OR uut_a_3_2 /= "000001100111010000101001010" OR uut_a_3_3 /= "000000000011010100000100010" OR uut_a_3_4 /= "111111110110000011110011010" OR uut_a_3_5 /= "000011100010111110100011001" OR uut_a_4_0 /= "111111111111111101101111010" OR uut_a_4_1 /= "000000000000000110110010001" OR uut_a_4_2 /= "111111111101100101000111000" OR uut_a_4_3 /= "111111111111111011000001111" OR uut_a_4_4 /= "000000000000001110111010010" OR uut_a_4_5 /= "111111111010101011100010001" OR uut_a_5_0 /= "000000000000110011101000010" OR uut_a_5_1 /= "111111111101100101000111000" OR uut_a_5_2 /= "000000110111010000101010000" OR uut_a_5_3 /= "000000000001110001011111010" OR uut_a_5_4 /= "111111111010101011100010001" OR uut_a_5_5 /= "000001111001011101111110010" THEN
              FAIL <= '1';
              FAIL_NUM <= "00110011";
              state <= "11111101";
            ELSE
              state <= "01000001";
            END IF;
            uut_rst <= '0';
          WHEN "01000001" =>
            uut_coord_shift <= "1000";
            uut_x <= "111101110001";
            uut_y <= "000000111011";
            uut_fx <= "0011111000";
            uut_fy <= "1110110011";
            uut_ft <= "1110111000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000001001011000010" OR uut_a_0_1 /= "000000000110011100101011000" OR uut_a_0_2 /= "111111111101010111001011100" OR uut_a_0_3 /= "111111111111101010100100000" OR uut_a_0_4 /= "111111110001010000110000000" OR uut_a_0_5 /= "000000000110000001111000000" OR uut_a_1_0 /= "000000000000000011001110010" OR uut_a_1_1 /= "000000000010001101110110110" OR uut_a_1_2 /= "111111111111000101111101111" OR uut_a_1_3 /= "111111111111111000101000011" OR uut_a_1_4 /= "111111111010111011110000100" OR uut_a_1_5 /= "000000000010000100101001010" OR uut_a_2_0 /= "111111111111111110101011100" OR uut_a_2_1 /= "111111111111000101111101111" OR uut_a_2_2 /= "000000000000010111101111011" OR uut_a_2_3 /= "000000000000000011000000111" OR uut_a_2_4 /= "000000000010000100101001010" OR uut_a_2_5 /= "111111111111001001101111001" OR uut_a_3_0 /= "111111111111101010100100000" OR uut_a_3_1 /= "111111110001010000110000000" OR uut_a_3_2 /= "000000000110000001111000000" OR uut_a_3_3 /= "000000000000110001000000000" OR uut_a_3_4 /= "000000100001101100000000000" OR uut_a_3_5 /= "111111110010001110000000000" OR uut_a_4_0 /= "111111111111111000101000011" OR uut_a_4_1 /= "111111111010111011110000100" OR uut_a_4_2 /= "000000000010000100101001010" OR uut_a_4_3 /= "000000000000010000110110000" OR uut_a_4_4 /= "000000001011100101001000000" OR uut_a_4_5 /= "111111111011010000110100000" OR uut_a_5_0 /= "000000000000000011000000111" OR uut_a_5_1 /= "000000000010000100101001010" OR uut_a_5_2 /= "111111111111001001101111001" OR uut_a_5_3 /= "111111111111111001000111000" OR uut_a_5_4 /= "111111111011010000110100000" OR uut_a_5_5 /= "000000000001111100000010000" THEN
              FAIL <= '1';
              FAIL_NUM <= "00110100";
              state <= "11111101";
            ELSE
              state <= "01000010";
            END IF;
            uut_rst <= '0';
          WHEN "01000010" =>
            uut_coord_shift <= "1000";
            uut_x <= "111010000000";
            uut_y <= "111000011010";
            uut_fx <= "1100101001";
            uut_fy <= "1101000101";
            uut_ft <= "0010011101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000010011101110100010" OR uut_a_0_1 /= "111110001100000110101000010" OR uut_a_0_2 /= "000010101011011000001111011" OR uut_a_0_3 /= "111111111011010010100000000" OR uut_a_0_4 /= "000011011101011010100000000" OR uut_a_0_5 /= "111010111000100101110000000" OR uut_a_1_0 /= "111111111111000110000011010" OR uut_a_1_1 /= "000000101010100011100100001" OR uut_a_1_2 /= "111111000001000100100110010" OR uut_a_1_3 /= "000000000001101110101101010" OR uut_a_1_4 /= "111110101110101100110001010" OR uut_a_1_5 /= "000001111000001110001000111" OR uut_a_2_0 /= "000000000001010101101100000" OR uut_a_2_1 /= "111111000001000100100110010" OR uut_a_2_2 /= "000001011101000011011010010" OR uut_a_2_3 /= "111111111101011100010010111" OR uut_a_2_4 /= "000001111000001110001000111" OR uut_a_2_5 /= "111101001110001110011111110" OR uut_a_3_0 /= "111111111011010010100000000" OR uut_a_3_1 /= "000011011101011010100000000" OR uut_a_3_2 /= "111010111000100101110000000" OR uut_a_3_3 /= "000000001001000000000000000" OR uut_a_3_4 /= "111001011001000000000000000" OR uut_a_3_5 /= "001001110001100000000000000" OR uut_a_4_0 /= "000000000001101110101101010" OR uut_a_4_1 /= "111110101110101100110001010" OR uut_a_4_2 /= "000001111000001110001000111" OR uut_a_4_3 /= "111111111100101100100000000" OR uut_a_4_4 /= "000010011011010100100000000" OR uut_a_4_5 /= "111100011010010100110000000" OR uut_a_5_0 /= "111111111101011100010010111" OR uut_a_5_1 /= "000001111000001110001000111" OR uut_a_5_2 /= "111101001110001110011111110" OR uut_a_5_3 /= "000000000100111000110000000" OR uut_a_5_4 /= "111100011010010100110000000" OR uut_a_5_5 /= "000101010011101000001000000" THEN
              FAIL <= '1';
              FAIL_NUM <= "00110101";
              state <= "11111101";
            ELSE
              state <= "01000011";
            END IF;
            uut_rst <= '0';
          WHEN "01000011" =>
            uut_coord_shift <= "1000";
            uut_x <= "000111010011";
            uut_y <= "000110111110";
            uut_fx <= "1111010101";
            uut_fy <= "1011110110";
            uut_ft <= "0100001110";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000011000011000010" OR uut_a_0_1 /= "111111011000011000100110000" OR uut_a_0_2 /= "111111010000001100011100101" OR uut_a_0_3 /= "111111111111001110111011110" OR uut_a_0_4 /= "000001001111101110111010000" OR uut_a_0_5 /= "000001100000001101110101011" OR uut_a_1_0 /= "111111111111101100001100010" OR uut_a_1_1 /= "000000100000001100000001001" OR uut_a_1_2 /= "000000100110110101111000101" OR uut_a_1_3 /= "000000000000100111110111011" OR uut_a_1_4 /= "111110111111001101111000111" OR uut_a_1_5 /= "111110110001110100110000101" OR uut_a_2_0 /= "111111111111101000000110001" OR uut_a_2_1 /= "000000100110110101111000101" OR uut_a_2_2 /= "000000101110110111110010111" OR uut_a_2_3 /= "000000000000110000000110111" OR uut_a_2_4 /= "111110110001110100110000101" OR uut_a_2_5 /= "111110100001101010011011111" OR uut_a_3_0 /= "111111111111001110111011110" OR uut_a_3_1 /= "000001001111101110111010000" OR uut_a_3_2 /= "000001100000001101110101011" OR uut_a_3_3 /= "000000000001100010110000010" OR uut_a_3_4 /= "111101011111100001100110000" OR uut_a_3_5 /= "111100111110010110011000101" OR uut_a_4_0 /= "000000000000100111110111011" OR uut_a_4_1 /= "111110111111001101111000111" OR uut_a_4_2 /= "111110110001110100110000101" OR uut_a_4_3 /= "111111111110101111110000110" OR uut_a_4_4 /= "000010000010011000101101001" OR uut_a_4_5 /= "000010011101010101110011111" OR uut_a_5_0 /= "000000000000110000000110111" OR uut_a_5_1 /= "111110110001110100110000101" OR uut_a_5_2 /= "111110100001101010011011111" OR uut_a_5_3 /= "111111111110011111001011001" OR uut_a_5_4 /= "000010011101010101110011111" OR uut_a_5_5 /= "000010111101110111100011010" THEN
              FAIL <= '1';
              FAIL_NUM <= "00110110";
              state <= "11111101";
            ELSE
              state <= "01000100";
            END IF;
            uut_rst <= '0';
          WHEN "01000100" =>
            uut_coord_shift <= "1000";
            uut_x <= "000100001001";
            uut_y <= "000011110110";
            uut_fx <= "0011111010";
            uut_fy <= "1001101100";
            uut_ft <= "0010111010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001000111001100010" OR uut_a_0_1 /= "000000001000010101111011111" OR uut_a_0_2 /= "111110010000110000110111000" OR uut_a_0_3 /= "111111111100110110100011100" OR uut_a_0_4 /= "111111101000011001001010010" OR uut_a_0_5 /= "000100111010110000100010000" OR uut_a_1_0 /= "000000000000000100001010111" OR uut_a_1_1 /= "000000000000011111010010010" OR uut_a_1_2 /= "111111111001011110110111001" OR uut_a_1_3 /= "111111111111110100001100100" OR uut_a_1_4 /= "111111111110100111011110010" OR uut_a_1_5 /= "000000010010011100010101111" OR uut_a_2_0 /= "111111111111001000011000011" OR uut_a_2_1 /= "111111111001011110110111001" OR uut_a_2_2 /= "000001010110111001110101000" OR uut_a_2_3 /= "000000000010011101011000010" OR uut_a_2_4 /= "000000010010011100010101111" OR uut_a_2_5 /= "111100001010000110000101011" OR uut_a_3_0 /= "111111111100110110100011100" OR uut_a_3_1 /= "111111101000011001001010010" OR uut_a_3_2 /= "000100111010110000100010000" OR uut_a_3_3 /= "000000001000111010000001000" OR uut_a_3_4 /= "000001000010110011000111100" OR uut_a_3_5 /= "110010000101010110011100000" OR uut_a_4_0 /= "111111111111110100001100100" OR uut_a_4_1 /= "111111111110100111011110010" OR uut_a_4_2 /= "000000010010011100010101111" OR uut_a_4_3 /= "000000000000100001011001100" OR uut_a_4_4 /= "000000000011111010011111101" OR uut_a_4_5 /= "111111001011110100000100001" OR uut_a_5_0 /= "000000000010011101011000010" OR uut_a_5_1 /= "000000010010011100010101111" OR uut_a_5_2 /= "111100001010000110000101011" OR uut_a_5_3 /= "111111111001000010101011001" OR uut_a_5_4 /= "111111001011110100000100001" OR uut_a_5_5 /= "001010110111110100011110001" THEN
              FAIL <= '1';
              FAIL_NUM <= "00110111";
              state <= "11111101";
            ELSE
              state <= "01000101";
            END IF;
            uut_rst <= '0';
          WHEN "01000101" =>
            uut_coord_shift <= "1000";
            uut_x <= "111111011011";
            uut_y <= "111011011010";
            uut_fx <= "1001100101";
            uut_fy <= "0101001011";
            uut_ft <= "1010110011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000111000011100100000" OR uut_a_0_1 /= "110100101100110010110110000" OR uut_a_0_2 /= "110101111010011010000010000" OR uut_a_0_3 /= "000000000110011101000011000" OR uut_a_0_4 /= "110101101010011110101100100" OR uut_a_0_5 /= "110110110001011110001101100" OR uut_a_1_0 /= "111111111010010110011001011" OR uut_a_1_1 /= "001001000011001000010010010" OR uut_a_1_2 /= "001000000100111110101001111" OR uut_a_1_3 /= "111111111010110101001111010" OR uut_a_1_4 /= "001000010001101110111010110" OR uut_a_1_5 /= "000111011000111000100011101" OR uut_a_2_0 /= "111111111010111101001101000" OR uut_a_2_1 /= "001000000100111110101001111" OR uut_a_2_2 /= "000111001101011111111001000" OR uut_a_2_3 /= "111111111011011000101111000" OR uut_a_2_4 /= "000111011000111000100011101" OR uut_a_2_5 /= "000110100110001000101001110" OR uut_a_3_0 /= "000000000110011101000011000" OR uut_a_3_1 /= "110101101010011110101100100" OR uut_a_3_2 /= "110110110001011110001101100" OR uut_a_3_3 /= "000000000101111001110100010" OR uut_a_3_4 /= "110110100010111001110100011" OR uut_a_3_5 /= "110111100011110101110011001" OR uut_a_4_0 /= "111111111010110101001111010" OR uut_a_4_1 /= "001000010001101110111010110" OR uut_a_4_2 /= "000111011000111000100011101" OR uut_a_4_3 /= "111111111011010001011100111" OR uut_a_4_4 /= "000111100100100011001100110" OR uut_a_4_5 /= "000110110000100011001010110" OR uut_a_5_0 /= "111111111011011000101111000" OR uut_a_5_1 /= "000111011000111000100011101" OR uut_a_5_2 /= "000110100110001000101001110" OR uut_a_5_3 /= "111111111011110001111010111" OR uut_a_5_4 /= "000110110000100011001010110" OR uut_a_5_5 /= "000110000010001000010010101" THEN
              FAIL <= '1';
              FAIL_NUM <= "00111000";
              state <= "11111101";
            ELSE
              state <= "01000110";
            END IF;
            uut_rst <= '0';
          WHEN "01000110" =>
            uut_coord_shift <= "1000";
            uut_x <= "111010101000";
            uut_y <= "000010101001";
            uut_fx <= "0110010100";
            uut_fy <= "0000010001";
            uut_ft <= "0011010000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000011111110000000010" OR uut_a_0_1 /= "111101000111011100110100011" OR uut_a_0_2 /= "111011100010001111101110000" OR uut_a_0_3 /= "111111111001101111100100100" OR uut_a_0_4 /= "000100100010111011111110110" OR uut_a_0_5 /= "000111000010011110111100000" OR uut_a_1_0 /= "111111111110100011101110011" OR uut_a_1_1 /= "000001000011000010110001111" OR uut_a_1_2 /= "000001100111110011110010100" OR uut_a_1_3 /= "000000000010010001011101111" OR uut_a_1_4 /= "111110010110010011101101011" OR uut_a_1_5 /= "111101011100010110010000101" OR uut_a_2_0 /= "111111111101110001000111110" OR uut_a_2_1 /= "000001100111110011110010100" OR uut_a_2_2 /= "000010100000101111001010001" OR uut_a_2_3 /= "000000000011100001001111011" OR uut_a_2_4 /= "111101011100010110010000101" OR uut_a_2_5 /= "111100000010100110100110010" OR uut_a_3_0 /= "111111111001101111100100100" OR uut_a_3_1 /= "000100100010111011111110110" OR uut_a_3_2 /= "000111000010011110111100000" OR uut_a_3_3 /= "000000001001110111010001000" OR uut_a_3_4 /= "111000110101010110001001100" OR uut_a_3_5 /= "110100111001110100111000000" OR uut_a_4_0 /= "000000000010010001011101111" OR uut_a_4_1 /= "111110010110010011101101011" OR uut_a_4_2 /= "111101011100010110010000101" OR uut_a_4_3 /= "111111111100011010101011000" OR uut_a_4_4 /= "000010100110100111101101000" OR uut_a_4_5 /= "000100000001111111100010101" OR uut_a_5_0 /= "000000000011100001001111011" OR uut_a_5_1 /= "111101011100010110010000101" OR uut_a_5_2 /= "111100000010100110100110010" OR uut_a_5_3 /= "111111111010011100111010011" OR uut_a_5_4 /= "000100000001111111100010101" OR uut_a_5_5 /= "000110001111011110010000100" THEN
              FAIL <= '1';
              FAIL_NUM <= "00111001";
              state <= "11111101";
            ELSE
              state <= "01000111";
            END IF;
            uut_rst <= '0';
          WHEN "01000111" =>
            uut_coord_shift <= "1000";
            uut_x <= "111010011110";
            uut_y <= "000111010000";
            uut_fx <= "0000101010";
            uut_fy <= "0010111000";
            uut_ft <= "1000100101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000101010011111100010" OR uut_a_0_1 /= "000001001010010111001011100" OR uut_a_0_2 /= "111001010100011010101101111" OR uut_a_0_3 /= "000000000111110010111101110" OR uut_a_0_4 /= "000001101101001001100000100" OR uut_a_0_5 /= "110110001100011001010101001" OR uut_a_1_0 /= "000000000000100101001011100" OR uut_a_1_1 /= "000000001000001000100010010" OR uut_a_1_2 /= "111111010001001110111011000" OR uut_a_1_3 /= "000000000000110110100100110" OR uut_a_1_4 /= "000000001011111100000010100" OR uut_a_1_5 /= "111110111011010110110001010" OR uut_a_2_0 /= "111111111100101010001101010" OR uut_a_2_1 /= "111111010001001110111011000" OR uut_a_2_2 /= "000100001100111010001100101" OR uut_a_2_3 /= "111111111011000110001100101" OR uut_a_2_4 /= "111110111011010110110001010" OR uut_a_2_5 /= "000110001010101101000100011" OR uut_a_3_0 /= "000000000111110010111101110" OR uut_a_3_1 /= "000001101101001001100000100" OR uut_a_3_2 /= "110110001100011001010101001" OR uut_a_3_3 /= "000000001011011100011000010" OR uut_a_3_4 /= "000010100000001101010011100" OR uut_a_3_5 /= "110001100110110011011111111" OR uut_a_4_0 /= "000000000000110110100100110" OR uut_a_4_1 /= "000000001011111100000010100" OR uut_a_4_2 /= "111110111011010110110001010" OR uut_a_4_3 /= "000000000001010000000110101" OR uut_a_4_4 /= "000000010001100001011101001" OR uut_a_4_5 /= "111110011011001111101000011" OR uut_a_5_0 /= "111111111011000110001100101" OR uut_a_5_1 /= "111110111011010110110001010" OR uut_a_5_2 /= "000110001010101101000100011" OR uut_a_5_3 /= "111111111000110011011001101" OR uut_a_5_4 /= "111110011011001111101000011" OR uut_a_5_5 /= "001001000011010110000111001" THEN
              FAIL <= '1';
              FAIL_NUM <= "00111010";
              state <= "11111101";
            ELSE
              state <= "01001000";
            END IF;
            uut_rst <= '0';
          WHEN "01001000" =>
            uut_coord_shift <= "1000";
            uut_x <= "000100111100";
            uut_y <= "000011111110";
            uut_fx <= "1001111011";
            uut_fy <= "0000011010";
            uut_ft <= "1101001110";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000010001110100000010" OR uut_a_0_1 /= "000001110100111001011101001" OR uut_a_0_2 /= "000000100000010010010011101" OR uut_a_0_3 /= "000000000011111111001010100" OR uut_a_0_4 /= "000011010001010100000111010" OR uut_a_0_5 /= "000000111001110011111000010" OR uut_a_1_0 /= "000000000000111010011100101" OR uut_a_1_1 /= "000000101111111100100100001" OR uut_a_1_2 /= "000000001101001111100000100" OR uut_a_1_3 /= "000000000001101000101010000" OR uut_a_1_4 /= "000001010101110110011111111" OR uut_a_1_5 /= "000000010111101101100001110" OR uut_a_2_0 /= "000000000000010000001001001" OR uut_a_2_1 /= "000000001101001111100000100" OR uut_a_2_2 /= "000000000011101010000100101" OR uut_a_2_3 /= "000000000000011100111001111" OR uut_a_2_4 /= "000000010111101101100001110" OR uut_a_2_5 /= "000000000110100011001000000" OR uut_a_3_0 /= "000000000011111111001010100" OR uut_a_3_1 /= "000011010001010100000111010" OR uut_a_3_2 /= "000000111001110011111000010" OR uut_a_3_3 /= "000000000111001000111001000" OR uut_a_3_4 /= "000101110110110010110000100" OR uut_a_3_5 /= "000001100111100000111010100" OR uut_a_4_0 /= "000000000001101000101010000" OR uut_a_4_1 /= "000001010101110110011111111" OR uut_a_4_2 /= "000000010111101101100001110" OR uut_a_4_3 /= "000000000010111011011001011" OR uut_a_4_4 /= "000010011001101110010100011" OR uut_a_4_5 /= "000000101010011101001111111" OR uut_a_5_0 /= "000000000000011100111001111" OR uut_a_5_1 /= "000000010111101101100001110" OR uut_a_5_2 /= "000000000110100011001000000" OR uut_a_5_3 /= "000000000000110011110000011" OR uut_a_5_4 /= "000000101010011101001111111" OR uut_a_5_5 /= "000000001011101110011110101" THEN
              FAIL <= '1';
              FAIL_NUM <= "00111011";
              state <= "11111101";
            ELSE
              state <= "01001001";
            END IF;
            uut_rst <= '0';
          WHEN "01001001" =>
            uut_coord_shift <= "1000";
            uut_x <= "000000101111";
            uut_y <= "111110011001";
            uut_fx <= "1110101001";
            uut_fy <= "1010111001";
            uut_ft <= "1100000110";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001111000001000000" OR uut_a_0_1 /= "000111010100010011001100000" OR uut_a_0_2 /= "111011000011101110111100000" OR uut_a_0_3 /= "000000000000110011010110000" OR uut_a_0_4 /= "000011001000001010010001000" OR uut_a_0_5 /= "111101111000110100100101000" OR uut_a_1_0 /= "000000000001110101000100110" OR uut_a_1_1 /= "000111001000011010001100110" OR uut_a_1_2 /= "111011001011110000110111101" OR uut_a_1_3 /= "000000000000110010000010100" OR uut_a_1_4 /= "000011000011000101000000010" OR uut_a_1_5 /= "111101111100010000001111100" OR uut_a_2_0 /= "111111111110110000111011101" OR uut_a_2_1 /= "111011001011110000110111101" OR uut_a_2_2 /= "000011010000001010101110110" OR uut_a_2_3 /= "111111111111011110001101001" OR uut_a_2_4 /= "111101111100010000001111100" OR uut_a_2_5 /= "000001011000111110011001001" OR uut_a_3_0 /= "000000000000110011010110000" OR uut_a_3_1 /= "000011001000001010010001000" OR uut_a_3_2 /= "111101111000110100100101000" OR uut_a_3_3 /= "000000000000010101111100100" OR uut_a_3_4 /= "000001010101100011010110110" OR uut_a_3_5 /= "111111000110001110001101110" OR uut_a_4_0 /= "000000000000110010000010100" OR uut_a_4_1 /= "000011000011000101000000010" OR uut_a_4_2 /= "111101111100010000001111100" OR uut_a_4_3 /= "000000000000010101011000110" OR uut_a_4_4 /= "000001010011011000010101010" OR uut_a_4_5 /= "111111000111101100000110101" OR uut_a_5_0 /= "111111111111011110001101001" OR uut_a_5_1 /= "111101111100010000001111100" OR uut_a_5_2 /= "000001011000111110011001001" OR uut_a_5_3 /= "111111111111110001100011100" OR uut_a_5_4 /= "111111000111101100000110101" OR uut_a_5_5 /= "000000100110000001111001001" THEN
              FAIL <= '1';
              FAIL_NUM <= "00111100";
              state <= "11111101";
            ELSE
              state <= "01001010";
            END IF;
            uut_rst <= '0';
          WHEN "01001010" =>
            uut_coord_shift <= "1000";
            uut_x <= "111000010110";
            uut_y <= "000110110001";
            uut_fx <= "0010011101";
            uut_fy <= "0110111011";
            uut_ft <= "1010100111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000111011100101000100" OR uut_a_0_1 /= "001010111100000011011111000" OR uut_a_0_2 /= "111010001111010110101011010" OR uut_a_0_3 /= "111111111110011111100001000" OR uut_a_0_4 /= "111101110010010010011110000" OR uut_a_0_5 /= "000001001010100111111110100" OR uut_a_1_0 /= "000000000010101111000000110" OR uut_a_1_1 /= "000100000001000011010001111" OR uut_a_1_2 /= "111101111000101000110100111" OR uut_a_1_3 /= "111111111111011100100100100" OR uut_a_1_4 /= "111111001011111101110010000" OR uut_a_1_5 /= "000000011011011001101011011" OR uut_a_2_0 /= "111111111110100011110101101" OR uut_a_2_1 /= "111101111000101000110100111" OR uut_a_2_2 /= "000001000111010001111111011" OR uut_a_2_3 /= "000000000000010010101001111" OR uut_a_2_4 /= "000000011011011001101011011" OR uut_a_2_5 /= "111111110001100100100001010" OR uut_a_3_0 /= "111111111110011111100001000" OR uut_a_3_1 /= "111101110010010010011110000" OR uut_a_3_2 /= "000001001010100111111110100" OR uut_a_3_3 /= "000000000000010011100010000" OR uut_a_3_4 /= "000000011100101011111100000" OR uut_a_3_5 /= "111111110000111001001101000" OR uut_a_4_0 /= "111111111111011100100100100" OR uut_a_4_1 /= "111111001011111101110010000" OR uut_a_4_2 /= "000000011011011001101011011" OR uut_a_4_3 /= "000000000000000111001010111" OR uut_a_4_4 /= "000000001010100010001000100" OR uut_a_4_5 /= "111111111010011101000000010" OR uut_a_5_0 /= "000000000000010010101001111" OR uut_a_5_1 /= "000000011011011001101011011" OR uut_a_5_2 /= "111111110001100100100001010" OR uut_a_5_3 /= "111111111111111100001110010" OR uut_a_5_4 /= "111111111010011101000000010" OR uut_a_5_5 /= "000000000010111010111100000" THEN
              FAIL <= '1';
              FAIL_NUM <= "00111101";
              state <= "11111101";
            ELSE
              state <= "01001011";
            END IF;
            uut_rst <= '0';
          WHEN "01001011" =>
            uut_coord_shift <= "1000";
            uut_x <= "000110101111";
            uut_y <= "000100101101";
            uut_fx <= "0001001111";
            uut_fy <= "1111000011";
            uut_ft <= "1100001000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000011101011001011001" OR uut_a_0_1 /= "110101110111011011110100011" OR uut_a_0_2 /= "111100100001101011111110111" OR uut_a_0_3 /= "111111111101001101000101000" OR uut_a_0_4 /= "000111101101011011101101100" OR uut_a_0_5 /= "000010101001001000110001100" OR uut_a_1_0 /= "111111111101011101110110111" OR uut_a_1_1 /= "000110111111001001111100011" OR uut_a_1_2 /= "000010011001010001100011001" OR uut_a_1_3 /= "000000000001111011010110111" OR uut_a_1_4 /= "111010101011110011010001010" OR uut_a_1_5 /= "111110001011011000110100110" OR uut_a_2_0 /= "111111111111001000011010111" OR uut_a_2_1 /= "000010011001010001100011001" OR uut_a_2_2 /= "000000110100100010011110110" OR uut_a_2_3 /= "000000000000101010010010001" OR uut_a_2_4 /= "111110001011011000110100110" OR uut_a_2_5 /= "111111011000000001110011010" OR uut_a_3_0 /= "111111111101001101000101000" OR uut_a_3_1 /= "000111101101011011101101100" OR uut_a_3_2 /= "000010101001001000110001100" OR uut_a_3_3 /= "000000000010001000001000000" OR uut_a_3_4 /= "111010001000100101111100000" OR uut_a_3_5 /= "111101111111010100011100000" OR uut_a_4_0 /= "000000000001111011010110111" OR uut_a_4_1 /= "111010101011110011010001010" OR uut_a_4_2 /= "111110001011011000110100110" OR uut_a_4_3 /= "111111111110100010001001011" OR uut_a_4_4 /= "000100000010110100110110000" OR uut_a_4_5 /= "000001011000101110000010001" OR uut_a_5_0 /= "000000000000101010010010001" OR uut_a_5_1 /= "111110001011011000110100110" OR uut_a_5_2 /= "111111011000000001110011010" OR uut_a_5_3 /= "111111111111011111110101000" OR uut_a_5_4 /= "000001011000101110000010001" OR uut_a_5_5 /= "000000011110011010010010111" THEN
              FAIL <= '1';
              FAIL_NUM <= "00111110";
              state <= "11111101";
            ELSE
              state <= "01001100";
            END IF;
            uut_rst <= '0';
          WHEN "01001100" =>
            uut_coord_shift <= "1000";
            uut_x <= "000100000001";
            uut_y <= "111011101011";
            uut_fx <= "1001000010";
            uut_fy <= "0100010010";
            uut_ft <= "0010101111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001010110111101001" OR uut_a_0_1 /= "111110011000101111011010100" OR uut_a_0_2 /= "000010000000011001010000010" OR uut_a_0_3 /= "111111111111110011001110011" OR uut_a_0_4 /= "000000001111001010111011100" OR uut_a_0_5 /= "111111101101001000101110011" OR uut_a_1_0 /= "111111111111100110001011110" OR uut_a_1_1 /= "000000011110101001111011001" OR uut_a_1_2 /= "111111011001111000100000001" OR uut_a_1_3 /= "000000000000000011110010101" OR uut_a_1_4 /= "111111111011011111110000010" OR uut_a_1_5 /= "000000000101100110011010001" OR uut_a_2_0 /= "000000000000100000000110010" OR uut_a_2_1 /= "111111011001111000100000001" OR uut_a_2_2 /= "000000101111011001010100101" OR uut_a_2_3 /= "111111111111111011010010001" OR uut_a_2_4 /= "000000000101100110011010001" OR uut_a_2_5 /= "111111111001000010010110001" OR uut_a_3_0 /= "111111111111110011001110011" OR uut_a_3_1 /= "000000001111001010111011100" OR uut_a_3_2 /= "111111101101001000101110011" OR uut_a_3_3 /= "000000000000000001111000001" OR uut_a_3_4 /= "111111111101110001010110100" OR uut_a_3_5 /= "000000000010110001010111110" OR uut_a_4_0 /= "000000000000000011110010101" OR uut_a_4_1 /= "111111111011011111110000010" OR uut_a_4_2 /= "000000000101100110011010001" OR uut_a_4_3 /= "111111111111111111011100010" OR uut_a_4_4 /= "000000000000101010010110010" OR uut_a_4_5 /= "111111111111001011010101111" OR uut_a_5_0 /= "111111111111111011010010001" OR uut_a_5_1 /= "000000000101100110011010001" OR uut_a_5_2 /= "111111111001000010010110001" OR uut_a_5_3 /= "000000000000000000101100010" OR uut_a_5_4 /= "111111111111001011010101111" OR uut_a_5_5 /= "000000000001000001011110011" THEN
              FAIL <= '1';
              FAIL_NUM <= "00111111";
              state <= "11111101";
            ELSE
              state <= "01001101";
            END IF;
            uut_rst <= '0';
          WHEN "01001101" =>
            uut_coord_shift <= "1000";
            uut_x <= "000011011100";
            uut_y <= "000010010001";
            uut_fx <= "1110101101";
            uut_fy <= "1110010000";
            uut_ft <= "0101000100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001010010111000100" OR uut_a_0_1 /= "000001000000000110101100110" OR uut_a_0_2 /= "111110010011001101110110000" OR uut_a_0_3 /= "000000000000010011101101110" OR uut_a_0_4 /= "000000001111001111111000101" OR uut_a_0_5 /= "111111100110000111111101000" OR uut_a_1_0 /= "000000000000010000000001101" OR uut_a_1_1 /= "000000001100011001010010111" OR uut_a_1_2 /= "111111101010111101110011010" OR uut_a_1_3 /= "000000000000000011110011111" OR uut_a_1_4 /= "000000000010111100101100100" OR uut_a_1_5 /= "111111111010111111110010011" OR uut_a_2_0 /= "111111111111100100110011011" OR uut_a_2_1 /= "111111101010111101110011010" OR uut_a_2_2 /= "000000100011101100011101010" OR uut_a_2_3 /= "111111111111111001100001111" OR uut_a_2_4 /= "111111111010111111110010011" OR uut_a_2_5 /= "000000001000011111011000111" OR uut_a_3_0 /= "000000000000010011101101110" OR uut_a_3_1 /= "000000001111001111111000101" OR uut_a_3_2 /= "111111100110000111111101000" OR uut_a_3_3 /= "000000000000000100101100001" OR uut_a_3_4 /= "000000000011101000001000001" OR uut_a_3_5 /= "111111111001110110000101100" OR uut_a_4_0 /= "000000000000000011110011111" OR uut_a_4_1 /= "000000000010111100101100100" OR uut_a_4_2 /= "111111111010111111110010011" OR uut_a_4_3 /= "000000000000000000111010000" OR uut_a_4_4 /= "000000000000101100111000100" OR uut_a_4_5 /= "111111111110110011110101010" OR uut_a_5_0 /= "111111111111111001100001111" OR uut_a_5_1 /= "111111111010111111110010011" OR uut_a_5_2 /= "000000001000011111011000111" OR uut_a_5_3 /= "111111111111111110011101100" OR uut_a_5_4 /= "111111111110110011110101010" OR uut_a_5_5 /= "000000000010000001010000001" THEN
              FAIL <= '1';
              FAIL_NUM <= "01000000";
              state <= "11111101";
            ELSE
              state <= "01001110";
            END IF;
            uut_rst <= '0';
          WHEN "01001110" =>
            uut_coord_shift <= "1000";
            uut_x <= "111101000110";
            uut_y <= "000101000010";
            uut_fx <= "0100101000";
            uut_fy <= "0101101001";
            uut_ft <= "0000000110";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001111000001000000" OR uut_a_0_1 /= "111101111001110011000100000" OR uut_a_0_2 /= "000000110111010111101100000" OR uut_a_0_3 /= "111111111111011010101101000" OR uut_a_0_4 /= "000000101001101010101110100" OR uut_a_0_5 /= "111111101110110011101111100" OR uut_a_1_0 /= "111111111111011110011100110" OR uut_a_1_1 /= "000000100101011110110111010" OR uut_a_1_2 /= "111111110000100010010000100" OR uut_a_1_3 /= "000000000000001010011010101" OR uut_a_1_4 /= "111111110100010111001100010" OR uut_a_1_5 /= "000000000100110011010011000" OR uut_a_2_0 /= "000000000000001101110101111" OR uut_a_2_1 /= "111111110000100010010000100" OR uut_a_2_2 /= "000000000110011000010110101" OR uut_a_2_3 /= "111111111111111011101100111" OR uut_a_2_4 /= "000000000100110011010011000" OR uut_a_2_5 /= "111111111110000001001101100" OR uut_a_3_0 /= "111111111111011010101101000" OR uut_a_3_1 /= "000000101001101010101110100" OR uut_a_3_2 /= "111111101110110011101111100" OR uut_a_3_3 /= "000000000000001011100101001" OR uut_a_3_4 /= "111111110011000100000001100" OR uut_a_3_5 /= "000000000101010101100111001" OR uut_a_4_0 /= "000000000000001010011010101" OR uut_a_4_1 /= "111111110100010111001100010" OR uut_a_4_2 /= "000000000100110011010011000" OR uut_a_4_3 /= "111111111111111100110001000" OR uut_a_4_4 /= "000000000011100111010000000" OR uut_a_4_5 /= "111111111110100000100101101" OR uut_a_5_0 /= "111111111111111011101100111" OR uut_a_5_1 /= "000000000100110011010011000" OR uut_a_5_2 /= "111111111110000001001101100" OR uut_a_5_3 /= "000000000000000001010101011" OR uut_a_5_4 /= "111111111110100000100101101" OR uut_a_5_5 /= "000000000000100111010111011" THEN
              FAIL <= '1';
              FAIL_NUM <= "01000001";
              state <= "11111101";
            ELSE
              state <= "01001111";
            END IF;
            uut_rst <= '0';
          WHEN "01001111" =>
            uut_coord_shift <= "1000";
            uut_x <= "000010001010";
            uut_y <= "000111001101";
            uut_fx <= "1111000111";
            uut_fy <= "1000111101";
            uut_ft <= "0101111000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001011010010010001" OR uut_a_0_1 /= "111011110001001001101000000" OR uut_a_0_2 /= "111010101001001101001011101" OR uut_a_0_3 /= "000000000001001110100001101" OR uut_a_0_4 /= "111100010100011011001000000" OR uut_a_0_5 /= "111011010101110110010101001" OR uut_a_1_0 /= "111111111110111100010010011" OR uut_a_1_1 /= "000011001011001000110010000" OR uut_a_1_2 /= "000100000001000110000111010" OR uut_a_1_3 /= "111111111111000101000110110" OR uut_a_1_4 /= "000010110000101011101010000" OR uut_a_1_5 /= "000011011111100111010000001" OR uut_a_2_0 /= "111111111110101010010011010" OR uut_a_2_1 /= "000100000001000110000111010" OR uut_a_2_2 /= "000101000101011000101111001" OR uut_a_2_3 /= "111111111110110101011101100" OR uut_a_2_4 /= "000011011111100111010000001" OR uut_a_2_5 /= "000100011011000000101011011" OR uut_a_3_0 /= "000000000001001110100001101" OR uut_a_3_1 /= "111100010100011011001000000" OR uut_a_3_2 /= "111011010101110110010101001" OR uut_a_3_3 /= "000000000001000100010011001" OR uut_a_3_4 /= "111100110011000110101000000" OR uut_a_3_5 /= "111011111100101011011000101" OR uut_a_4_0 /= "111111111111000101000110110" OR uut_a_4_1 /= "000010110000101011101010000" OR uut_a_4_2 /= "000011011111100111010000001" OR uut_a_4_3 /= "111111111111001100110001101" OR uut_a_4_4 /= "000010011001101011000010000" OR uut_a_4_5 /= "000011000010011111011101100" OR uut_a_5_0 /= "111111111110110101011101100" OR uut_a_5_1 /= "000011011111100111010000001" OR uut_a_5_2 /= "000100011011000000101011011" OR uut_a_5_3 /= "111111111110111111001010110" OR uut_a_5_4 /= "000011000010011111011101100" OR uut_a_5_5 /= "000011110110001001110100011" THEN
              FAIL <= '1';
              FAIL_NUM <= "01000010";
              state <= "11111101";
            ELSE
              state <= "01010000";
            END IF;
            uut_rst <= '0';
          WHEN "01010000" =>
            uut_coord_shift <= "1001";
            uut_x <= "000100001100";
            uut_y <= "111011011000";
            uut_fx <= "0111111101";
            uut_fy <= "1011100110";
            uut_ft <= "0010011100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000011100111001" OR uut_a_0_1 /= "000000001101001011001111101" OR uut_a_0_2 /= "000000001100100101010100111" OR uut_a_0_3 /= "000000000000010110010101110" OR uut_a_0_4 /= "000001010001100000010110101" OR uut_a_0_5 /= "000001001101110101110010010" OR uut_a_1_0 /= "000000000000000011010010110" OR uut_a_1_1 /= "000000001100000001001000011" OR uut_a_1_2 /= "000000001011011110100010111" OR uut_a_1_3 /= "000000000000010100011000000" OR uut_a_1_4 /= "000001001010010101111000101" OR uut_a_1_5 /= "000001000110111111111011101" OR uut_a_2_0 /= "000000000000000011001001010" OR uut_a_2_1 /= "000000001011011110100010111" OR uut_a_2_2 /= "000000001010111101100000111" OR uut_a_2_3 /= "000000000000010011011101011" OR uut_a_2_4 /= "000001000110111111111011101" OR uut_a_2_5 /= "000001000011110011100110100" OR uut_a_3_0 /= "000000000000010110010101110" OR uut_a_3_1 /= "000001010001100000010110101" OR uut_a_3_2 /= "000001001101110101110010010" OR uut_a_3_3 /= "000000000010001010001100100" OR uut_a_3_4 /= "000111111000001100100110110" OR uut_a_3_5 /= "000111100001100001100011100" OR uut_a_4_0 /= "000000000000010100011000000" OR uut_a_4_1 /= "000001001010010101111000101" OR uut_a_4_2 /= "000001000110111111111011101" OR uut_a_4_3 /= "000000000001111110000011001" OR uut_a_4_4 /= "000111001011111000011111110" OR uut_a_4_5 /= "000110110111001100111110110" OR uut_a_5_0 /= "000000000000010011011101011" OR uut_a_5_1 /= "000001000110111111111011101" OR uut_a_5_2 /= "000001000011110011100110100" OR uut_a_5_3 /= "000000000001111000011000011" OR uut_a_5_4 /= "000110110111001100111110110" OR uut_a_5_5 /= "000110100011011100111110101" THEN
              FAIL <= '1';
              FAIL_NUM <= "01000011";
              state <= "11111101";
            ELSE
              state <= "01010001";
            END IF;
            uut_rst <= '0';
          WHEN "01010001" =>
            uut_coord_shift <= "1001";
            uut_x <= "000011010111";
            uut_y <= "111100011010";
            uut_fx <= "1010010010";
            uut_fy <= "1000011010";
            uut_ft <= "1110101111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001111010000100100" OR uut_a_0_1 /= "000011111100101110010100010" OR uut_a_0_2 /= "000011101010100110101001100" OR uut_a_0_3 /= "111111111100111010101111000" OR uut_a_0_4 /= "111001100111100110010011100" OR uut_a_0_5 /= "111010000100111000010101000" OR uut_a_1_0 /= "000000000000111111001011100" OR uut_a_1_1 /= "000010000010110011011110001" OR uut_a_1_2 /= "000001111001011011010000001" OR uut_a_1_3 /= "111111111110011001111001100" OR uut_a_1_4 /= "111100101100100111101100110" OR uut_a_1_5 /= "111100111011110001101001110" OR uut_a_2_0 /= "000000000000111010101001101" OR uut_a_2_1 /= "000001111001011011010000001" OR uut_a_2_2 /= "000001110000101110000100011" OR uut_a_2_3 /= "111111111110100001001110000" OR uut_a_2_4 /= "111100111011110001101001110" OR uut_a_2_5 /= "111101001001110110000100000" OR uut_a_3_0 /= "111111111100111010101111000" OR uut_a_3_1 /= "111001100111100110010011100" OR uut_a_3_2 /= "111010000100111000010101000" OR uut_a_3_3 /= "000000000100111110110010000" OR uut_a_3_4 /= "001010010011111110100001000" OR uut_a_3_5 /= "001001100100101010000110000" OR uut_a_4_0 /= "111111111110011001111001100" OR uut_a_4_1 /= "111100101100100111101100110" OR uut_a_4_2 /= "111100111011110001101001110" OR uut_a_4_3 /= "000000000010100100111111101" OR uut_a_4_4 /= "000101010101100101101110110" OR uut_a_4_5 /= "000100111101000110010010010" OR uut_a_5_0 /= "111111111110100001001110000" OR uut_a_5_1 /= "111100111011110001101001110" OR uut_a_5_2 /= "111101001001110110000100000" OR uut_a_5_3 /= "000000000010011001001010100" OR uut_a_5_4 /= "000100111101000110010010010" OR uut_a_5_5 /= "000100100110010111001110011" THEN
              FAIL <= '1';
              FAIL_NUM <= "01000100";
              state <= "11111101";
            ELSE
              state <= "01010010";
            END IF;
            uut_rst <= '0';
          WHEN "01010010" =>
            uut_coord_shift <= "1001";
            uut_x <= "110101111010";
            uut_y <= "000111001110";
            uut_fx <= "1101111011";
            uut_fy <= "0101011110";
            uut_ft <= "0011110000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000101001001111011001" OR uut_a_0_1 /= "111110100000101000011010001" OR uut_a_0_2 /= "110100001010001101001100101" OR uut_a_0_3 /= "111111111011110110010010111" OR uut_a_0_4 /= "000001001100110011100010110" OR uut_a_0_5 /= "001001100010010010101001011" OR uut_a_1_0 /= "111111111111101000001010000" OR uut_a_1_1 /= "000000000110111001000101000" OR uut_a_1_2 /= "000000110110110000110010111" OR uut_a_1_3 /= "000000000000010011001100111" OR uut_a_1_4 /= "111111111010011100110001100" OR uut_a_1_5 /= "111111010011111001011001110" OR uut_a_2_0 /= "111111111101000010100011010" OR uut_a_2_1 /= "000000110110110000110010111" OR uut_a_2_2 /= "000110110011001000111011000" OR uut_a_2_3 /= "000000000010011000100100101" OR uut_a_2_4 /= "111111010011111001011001110" OR uut_a_2_5 /= "111010100001100011110010101" OR uut_a_3_0 /= "111111111011110110010010111" OR uut_a_3_1 /= "000001001100110011100010110" OR uut_a_3_2 /= "001001100010010010101001011" OR uut_a_3_3 /= "000000000011010101111111001" OR uut_a_3_4 /= "111111000010001001010000001" OR uut_a_3_5 /= "111000010100100000000000101" OR uut_a_4_0 /= "000000000000010011001100111" OR uut_a_4_1 /= "111111111010011100110001100" OR uut_a_4_2 /= "111111010011111001011001110" OR uut_a_4_3 /= "111111111111110000100010010" OR uut_a_4_4 /= "000000000100011110000101001" OR uut_a_4_5 /= "000000100011100001001011111" OR uut_a_5_0 /= "000000000010011000100100101" OR uut_a_5_1 /= "111111010011111001011001110" OR uut_a_5_2 /= "111010100001100011110010101" OR uut_a_5_3 /= "111111111110000101001000000" OR uut_a_5_4 /= "000000100011100001001011111" OR uut_a_5_5 /= "000100011010001110100111101" THEN
              FAIL <= '1';
              FAIL_NUM <= "01000101";
              state <= "11111101";
            ELSE
              state <= "01010011";
            END IF;
            uut_rst <= '0';
          WHEN "01010011" =>
            uut_coord_shift <= "1001";
            uut_x <= "000010010001";
            uut_y <= "110101101011";
            uut_fx <= "0111010100";
            uut_fy <= "1100010000";
            uut_ft <= "0110110011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000100111110110010000" OR uut_a_0_1 /= "110010100111010001101000000" OR uut_a_0_2 /= "000110100100111001000001000" OR uut_a_0_3 /= "000000000000001101011010100" OR uut_a_0_4 /= "111111011011111100110010000" OR uut_a_0_5 /= "000000010001101101011111010" OR uut_a_1_0 /= "111111111100101001110100011" OR uut_a_1_1 /= "001000111111100111001010001" OR uut_a_1_2 /= "111011100101001101101100010" OR uut_a_1_3 /= "111111111111110110111111001" OR uut_a_1_4 /= "000000011000001110001010011" OR uut_a_1_5 /= "111111110100000110011100000" OR uut_a_2_0 /= "000000000001101001001110010" OR uut_a_2_1 /= "111011100101001101101100010" OR uut_a_2_2 /= "000010001010111011010100011" OR uut_a_2_3 /= "000000000000000100011011010" OR uut_a_2_4 /= "111111110100000110011100000" OR uut_a_2_5 /= "000000000101110110001000111" OR uut_a_3_0 /= "000000000000001101011010100" OR uut_a_3_1 /= "111111011011111100110010000" OR uut_a_3_2 /= "000000010001101101011111010" OR uut_a_3_3 /= "000000000000000000100100001" OR uut_a_3_4 /= "111111111110011110111010100" OR uut_a_3_5 /= "000000000000101111101100100" OR uut_a_4_0 /= "111111111111110110111111001" OR uut_a_4_1 /= "000000011000001110001010011" OR uut_a_4_2 /= "111111110100000110011100000" OR uut_a_4_3 /= "111111111111111111100111101" OR uut_a_4_4 /= "000000000001000001001110101" OR uut_a_4_5 /= "111111111111011111111101000" OR uut_a_5_0 /= "000000000000000100011011010" OR uut_a_5_1 /= "111111110100000110011100000" OR uut_a_5_2 /= "000000000101110110001000111" OR uut_a_5_3 /= "000000000000000000001011111" OR uut_a_5_4 /= "111111111111011111111101000" OR uut_a_5_5 /= "000000000000001111101111100" THEN
              FAIL <= '1';
              FAIL_NUM <= "01000110";
              state <= "11111101";
            ELSE
              state <= "01010100";
            END IF;
            uut_rst <= '0';
          WHEN "01010100" =>
            uut_coord_shift <= "1001";
            uut_x <= "110111001011";
            uut_y <= "111011111110";
            uut_fx <= "1001011010";
            uut_fy <= "0010001111";
            uut_ft <= "1010111001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000011011100100" OR uut_a_0_1 /= "111111110110011110001011100" OR uut_a_0_2 /= "000000001100011111010100000" OR uut_a_0_3 /= "000000000000001111000110000" OR uut_a_0_4 /= "111111010110010000011010000" OR uut_a_0_5 /= "000000110110101101110000000" OR uut_a_1_0 /= "111111111111111101100111100" OR uut_a_1_1 /= "000000000110100101101000100" OR uut_a_1_2 /= "111111110111010111010110011" OR uut_a_1_3 /= "111111111111110101100100000" OR uut_a_1_4 /= "000000011100110111001010000" OR uut_a_1_5 /= "111111011010001010110111100" OR uut_a_2_0 /= "000000000000000011000111110" OR uut_a_2_1 /= "111111110111010111010110011" OR uut_a_2_2 /= "000000001011010100011000001" OR uut_a_2_3 /= "000000000000001101101011011" OR uut_a_2_4 /= "111111011010001010110111100" OR uut_a_2_5 /= "000000110001100101011101100" OR uut_a_3_0 /= "000000000000001111000110000" OR uut_a_3_1 /= "111111010110010000011010000" OR uut_a_3_2 /= "000000110110101101110000000" OR uut_a_3_3 /= "000000000001000010001000000" OR uut_a_3_4 /= "111101001001000111111000000" OR uut_a_3_5 /= "000011101111101101000000000" OR uut_a_4_0 /= "111111111111110101100100000" OR uut_a_4_1 /= "000000011100110111001010000" OR uut_a_4_2 /= "111111011010001010110111100" OR uut_a_4_3 /= "111111111111010010010001111" OR uut_a_4_4 /= "000001111110011100010011100" OR uut_a_4_5 /= "111101011010010001001000110" OR uut_a_5_0 /= "000000000000001101101011011" OR uut_a_5_1 /= "111111011010001010110111100" OR uut_a_5_2 /= "000000110001100101011101100" OR uut_a_5_3 /= "000000000000111011111011010" OR uut_a_5_4 /= "111101011010010001001000110" OR uut_a_5_5 /= "000011011001001110110010000" THEN
              FAIL <= '1';
              FAIL_NUM <= "01000111";
              state <= "11111101";
            ELSE
              state <= "01010101";
            END IF;
            uut_rst <= '0';
          WHEN "01010101" =>
            uut_coord_shift <= "1001";
            uut_x <= "110001011101";
            uut_y <= "000111001001";
            uut_fx <= "1101100100";
            uut_fy <= "0010100100";
            uut_ft <= "1110001001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000100100111100011001" OR uut_a_0_1 /= "001011011001101000101101110" OR uut_a_0_2 /= "001001001010011110101100111" OR uut_a_0_3 /= "111111111111101100001111110" OR uut_a_0_4 /= "111111001111001110111000100" OR uut_a_0_5 /= "111111011000110011010000010" OR uut_a_1_0 /= "000000000010110110011010001" OR uut_a_1_1 /= "000111000010010100101000001" OR uut_a_1_2 /= "000101101001111101111100101" OR uut_a_1_3 /= "111111111111110011110011101" OR uut_a_1_4 /= "111111100001111001101011110" OR uut_a_1_5 /= "111111100111110011101000100" OR uut_a_2_0 /= "000000000010010010100111101" OR uut_a_2_1 /= "000101101001111101111100101" OR uut_a_2_2 /= "000100100010111100101110110" OR uut_a_2_3 /= "111111111111110110001100110" OR uut_a_2_4 /= "111111100111110011101000100" OR uut_a_2_5 /= "111111101100100011011011010" OR uut_a_3_0 /= "111111111111101100001111110" OR uut_a_3_1 /= "111111001111001110111000100" OR uut_a_3_2 /= "111111011000110011010000010" OR uut_a_3_3 /= "000000000000000001010100100" OR uut_a_3_4 /= "000000000011010000100111000" OR uut_a_3_5 /= "000000000010100111101011100" OR uut_a_4_0 /= "111111111111110011110011101" OR uut_a_4_1 /= "111111100001111001101011110" OR uut_a_4_2 /= "111111100111110011101000100" OR uut_a_4_3 /= "000000000000000000110100001" OR uut_a_4_4 /= "000000000010000000110000000" OR uut_a_4_5 /= "000000000001100111011111010" OR uut_a_5_0 /= "111111111111110110001100110" OR uut_a_5_1 /= "111111100111110011101000100" OR uut_a_5_2 /= "111111101100100011011011010" OR uut_a_5_3 /= "000000000000000000101001111" OR uut_a_5_4 /= "000000000001100111011111010" OR uut_a_5_5 /= "000000000001010011001011110" THEN
              FAIL <= '1';
              FAIL_NUM <= "01001000";
              state <= "11111101";
            ELSE
              state <= "01010110";
            END IF;
            uut_rst <= '0';
          WHEN "01010110" =>
            uut_coord_shift <= "1001";
            uut_x <= "000100000100";
            uut_y <= "110000101101";
            uut_fx <= "0110100100";
            uut_fy <= "0100110100";
            uut_ft <= "0011111100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000001110110010001" OR uut_a_0_1 /= "000000000101011011011001111" OR uut_a_0_2 /= "111111110100000110101010100" OR uut_a_0_3 /= "000000000000110111100100001" OR uut_a_0_4 /= "000000010100011001110000111" OR uut_a_0_5 /= "111111010011010010011011100" OR uut_a_1_0 /= "000000000000000001010110110" OR uut_a_1_1 /= "000000000000011111111001000" OR uut_a_1_2 /= "111111111110111010000111001" OR uut_a_1_3 /= "000000000000000101000110011" OR uut_a_1_4 /= "000000000001110111110111010" OR uut_a_1_5 /= "111111111011111001010100010" OR uut_a_2_0 /= "111111111111111101000001101" OR uut_a_2_1 /= "111111111110111010000111001" OR uut_a_2_2 /= "000000000010011001001010001" OR uut_a_2_3 /= "111111111111110100110100100" OR uut_a_2_4 /= "111111111011111001010100010" OR uut_a_2_5 /= "000000001000111111101010101" OR uut_a_3_0 /= "000000000000110111100100001" OR uut_a_3_1 /= "000000010100011001110000111" OR uut_a_3_2 /= "111111010011010010011011100" OR uut_a_3_3 /= "000000000011010000110110001" OR uut_a_3_4 /= "000001001100101011110111111" OR uut_a_3_5 /= "111101010111111100011100100" OR uut_a_4_0 /= "000000000000000101000110011" OR uut_a_4_1 /= "000000000001110111110111010" OR uut_a_4_2 /= "111111111011111001010100010" OR uut_a_4_3 /= "000000000000010011001010111" OR uut_a_4_4 /= "000000000111000010100001110" OR uut_a_4_5 /= "111111110000100100101011000" OR uut_a_5_0 /= "111111111111110100110100100" OR uut_a_5_1 /= "111111111011111001010100010" OR uut_a_5_2 /= "000000001000111111101010101" OR uut_a_5_3 /= "111111111111010101111111000" OR uut_a_5_4 /= "111111110000100100101011000" OR uut_a_5_5 /= "000000100001110011101101110" THEN
              FAIL <= '1';
              FAIL_NUM <= "01001001";
              state <= "11111101";
            ELSE
              state <= "01010111";
            END IF;
            uut_rst <= '0';
          WHEN "01010111" =>
            uut_coord_shift <= "1001";
            uut_x <= "001010000001";
            uut_y <= "111100010010";
            uut_fx <= "0001111000";
            uut_fy <= "0001001101";
            uut_ft <= "0000011111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000110000001001001" OR uut_a_0_1 /= "111101000111101101000100011" OR uut_a_0_2 /= "000010100010110110110111100" OR uut_a_0_3 /= "000000000010000111110101111" OR uut_a_0_4 /= "110111110111111110110000101" OR uut_a_0_5 /= "000111001011100001101111111" OR uut_a_1_0 /= "111111111111010001111011010" OR uut_a_1_1 /= "000010110000011000000111100" OR uut_a_1_2 /= "111101100100001000111111010" OR uut_a_1_3 /= "111111111101111101111111101" OR uut_a_1_4 /= "000111110001101011001011111" OR uut_a_1_5 /= "111001001000001101111100110" OR uut_a_2_0 /= "000000000000101000101101101" OR uut_a_2_1 /= "111101100100001000111111010" OR uut_a_2_2 /= "000010001001101110101001101" OR uut_a_2_3 /= "000000000001110010111000011" OR uut_a_2_4 /= "111001001000001101111100110" OR uut_a_2_5 /= "000110000100100111111010101" OR uut_a_3_0 /= "000000000010000111110101111" OR uut_a_3_1 /= "110111110111111110110000101" OR uut_a_3_2 /= "000111001011100001101111111" OR uut_a_3_3 /= "000000000101111111010011001" OR uut_a_3_4 /= "101001000100101011110010011" OR uut_a_3_5 /= "010100010000101000001100100" OR uut_a_4_0 /= "111111111101111101111111101" OR uut_a_4_1 /= "000111110001101011001011111" OR uut_a_4_2 /= "111001001000001101111100110" OR uut_a_4_3 /= "111111111010010001001010111" OR uut_a_4_4 /= "010101111100010001000110000" OR uut_a_4_5 /= "101100100111000101100001111" OR uut_a_5_0 /= "000000000001110010111000011" OR uut_a_5_1 /= "111001001000001101111100110" OR uut_a_5_2 /= "000110000100100111111010101" OR uut_a_5_3 /= "000000000101000100001010000" OR uut_a_5_4 /= "101100100111000101100001111" OR uut_a_5_5 /= "010001001000100011111111100" THEN
              FAIL <= '1';
              FAIL_NUM <= "01001010";
              state <= "11111101";
            ELSE
              state <= "01011000";
            END IF;
            uut_rst <= '0';
          WHEN "01011000" =>
            uut_coord_shift <= "1001";
            uut_x <= "111000110100";
            uut_y <= "110111111110";
            uut_fx <= "1111001110";
            uut_fy <= "1011101001";
            uut_ft <= "0100111000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000001100001100001" OR uut_a_0_1 /= "000000101001000010110100111" OR uut_a_0_2 /= "000000011100101010100000110" OR uut_a_0_3 /= "111111111111110110100101101" OR uut_a_0_4 /= "111111100000010011101100001" OR uut_a_0_5 /= "111111101001110111011110100" OR uut_a_1_0 /= "000000000000001010010000101" OR uut_a_1_1 /= "000000100010100011010000010" OR uut_a_1_2 /= "000000011000001000010010010" OR uut_a_1_3 /= "111111111111111000000100111" OR uut_a_1_4 /= "111111100101010100100100110" OR uut_a_1_5 /= "111111101101010111100100110" OR uut_a_2_0 /= "000000000000000111001010101" OR uut_a_2_1 /= "000000011000001000010010010" OR uut_a_2_2 /= "000000010000110110011111100" OR uut_a_2_3 /= "111111111111111010011101110" OR uut_a_2_4 /= "111111101101010111100100110" OR uut_a_2_5 /= "111111110010111111001111010" OR uut_a_3_0 /= "111111111111110110100101101" OR uut_a_3_1 /= "111111100000010011101100001" OR uut_a_3_2 /= "111111101001110111011110100" OR uut_a_3_3 /= "000000000000000111010001001" OR uut_a_3_4 /= "000000011000011110001010011" OR uut_a_3_5 /= "000000010001000101110001010" OR uut_a_4_0 /= "111111111111111000000100111" OR uut_a_4_1 /= "111111100101010100100100110" OR uut_a_4_2 /= "111111101101010111100100110" OR uut_a_4_3 /= "000000000000000110000111100" OR uut_a_4_4 /= "000000010100100110011001000" OR uut_a_4_5 /= "000000001110011000101110111" OR uut_a_5_0 /= "111111111111111010011101110" OR uut_a_5_1 /= "111111101101010111100100110" OR uut_a_5_2 /= "111111110010111111001111010" OR uut_a_5_3 /= "000000000000000100010001011" OR uut_a_5_4 /= "000000001110011000101110111" OR uut_a_5_5 /= "000000001010000011000001000" THEN
              FAIL <= '1';
              FAIL_NUM <= "01001011";
              state <= "11111101";
            ELSE
              state <= "01011001";
            END IF;
            uut_rst <= '0';
          WHEN "01011001" =>
            uut_coord_shift <= "1001";
            uut_x <= "001111100011";
            uut_y <= "110000111110";
            uut_fx <= "0000100101";
            uut_fy <= "1001011001";
            uut_ft <= "0100110101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000110000100100000100" OR uut_a_0_1 /= "001100001100000011010000010" OR uut_a_0_2 /= "110010110111001111101010110" OR uut_a_0_3 /= "111111111100010001010100100" OR uut_a_0_4 /= "111000100000110001101010010" OR uut_a_0_5 /= "001000000100100001001000110" OR uut_a_1_0 /= "000000000011000011000000110" OR uut_a_1_1 /= "000110000111100011001000100" OR uut_a_1_2 /= "111001011001111110101111010" OR uut_a_1_3 /= "111111111110001000001100011" OR uut_a_1_4 /= "111100001111011100111011010" OR uut_a_1_5 /= "000100000011010001001000100" OR uut_a_2_0 /= "111111111100101101110011111" OR uut_a_2_1 /= "111001011001111110101111010" OR uut_a_2_2 /= "000111000110110111001001011" OR uut_a_2_3 /= "000000000010000001001000010" OR uut_a_2_4 /= "000100000011010001001000100" OR uut_a_2_5 /= "111011101000100011100100101" OR uut_a_3_0 /= "111111111100010001010100100" OR uut_a_3_1 /= "111000100000110001101010010" OR uut_a_3_2 /= "001000000100100001001000110" OR uut_a_3_3 /= "000000000010010010101000100" OR uut_a_3_4 /= "000100100110011010010100010" OR uut_a_3_5 /= "111011000010101011010110110" OR uut_a_4_0 /= "111111111110001000001100011" OR uut_a_4_1 /= "111100001111011100111011010" OR uut_a_4_2 /= "000100000011010001001000100" OR uut_a_4_3 /= "000000000001001001100110100" OR uut_a_4_4 /= "000010010011110001111101011" OR uut_a_4_5 /= "111101100000101110000000110" OR uut_a_5_0 /= "000000000010000001001000010" OR uut_a_5_1 /= "000100000011010001001000100" OR uut_a_5_2 /= "111011101000100011100100101" OR uut_a_5_3 /= "111111111110110000101010110" OR uut_a_5_4 /= "111101100000101110000000110" OR uut_a_5_5 /= "000010101011101011010010110" THEN
              FAIL <= '1';
              FAIL_NUM <= "01001100";
              state <= "11111101";
            ELSE
              state <= "01011010";
            END IF;
            uut_rst <= '0';
          WHEN "01011010" =>
            uut_coord_shift <= "1001";
            uut_x <= "001111101001";
            uut_y <= "110010001010";
            uut_fx <= "0111000010";
            uut_fy <= "1000010011";
            uut_ft <= "0010111100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000001101011101001" OR uut_a_0_1 /= "000000010111001000000011110" OR uut_a_0_2 /= "000000001111001111011111100" OR uut_a_0_3 /= "000000000000010010001010000" OR uut_a_0_4 /= "000000011111001101001100000" OR uut_a_0_5 /= "000000010100100100010101000" OR uut_a_1_0 /= "000000000000000101110010000" OR uut_a_1_1 /= "000000001001111011111101100" OR uut_a_1_2 /= "000000000110100011001010000" OR uut_a_1_3 /= "000000000000000111110011010" OR uut_a_1_4 /= "000000001101011010001010101" OR uut_a_1_5 /= "000000001000110101100111000" OR uut_a_2_0 /= "000000000000000011110011110" OR uut_a_2_1 /= "000000000110100011001010000" OR uut_a_2_2 /= "000000000100010100010000110" OR uut_a_2_3 /= "000000000000000101001001000" OR uut_a_2_4 /= "000000001000110101100111000" OR uut_a_2_5 /= "000000000101110100110010011" OR uut_a_3_0 /= "000000000000010010001010000" OR uut_a_3_1 /= "000000011111001101001100000" OR uut_a_3_2 /= "000000010100100100010101000" OR uut_a_3_3 /= "000000000000011000100000000" OR uut_a_3_4 /= "000000101010000111000000000" OR uut_a_3_5 /= "000000011011110000010000000" OR uut_a_4_0 /= "000000000000000111110011010" OR uut_a_4_1 /= "000000001101011010001010101" OR uut_a_4_2 /= "000000001000110101100111000" OR uut_a_4_3 /= "000000000000001010100001110" OR uut_a_4_4 /= "000000010010000110000000100" OR uut_a_4_5 /= "000000001011111011001110111" OR uut_a_5_0 /= "000000000000000101001001000" OR uut_a_5_1 /= "000000001000110101100111000" OR uut_a_5_2 /= "000000000101110100110010011" OR uut_a_5_3 /= "000000000000000110111100000" OR uut_a_5_4 /= "000000001011111011001110111" OR uut_a_5_5 /= "000000000111110111000010100" THEN
              FAIL <= '1';
              FAIL_NUM <= "01001101";
              state <= "11111101";
            ELSE
              state <= "01011011";
            END IF;
            uut_rst <= '0';
          WHEN "01011011" =>
            uut_coord_shift <= "1001";
            uut_x <= "001001000101";
            uut_y <= "000001000101";
            uut_fx <= "0110001011";
            uut_fy <= "0110011001";
            uut_ft <= "0010000001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000010101011001000000" OR uut_a_0_1 /= "111100000111010101011000000" OR uut_a_0_2 /= "000110101110011111001000000" OR uut_a_0_3 /= "000000000011010000101101000" OR uut_a_0_4 /= "111011010000101110100111000" OR uut_a_0_5 /= "001000001101000001001101000" OR uut_a_1_0 /= "111111111111000001110101010" OR uut_a_1_1 /= "000001011010010101011111000" OR uut_a_1_2 /= "111101100011100111001100010" OR uut_a_1_3 /= "111111111110110100001011101" OR uut_a_1_4 /= "000001101110001011000100010" OR uut_a_1_5 /= "111101000001010001010100000" OR uut_a_2_0 /= "000000000001101011100111110" OR uut_a_2_1 /= "111101100011100111001100010" OR uut_a_2_2 /= "000100001110101111000100110" OR uut_a_2_3 /= "000000000010000011010000010" OR uut_a_2_4 /= "111101000001010001010100000" OR uut_a_2_5 /= "000101001010001100000000011" OR uut_a_3_0 /= "000000000011010000101101000" OR uut_a_3_1 /= "111011010000101110100111000" OR uut_a_3_2 /= "001000001101000001001101000" OR uut_a_3_3 /= "000000000011111110100010001" OR uut_a_3_4 /= "111010001110001000011010011" OR uut_a_3_5 /= "001010000000010011110110001" OR uut_a_4_0 /= "111111111110110100001011101" OR uut_a_4_1 /= "000001101110001011000100010" OR uut_a_4_2 /= "111101000001010001010100000" OR uut_a_4_3 /= "111111111110100011100010000" OR uut_a_4_4 /= "000010000110010111011100011" OR uut_a_4_5 /= "111100010111011000110010100" OR uut_a_5_0 /= "000000000010000011010000010" OR uut_a_5_1 /= "111101000001010001010100000" OR uut_a_5_2 /= "000101001010001100000000011" OR uut_a_5_3 /= "000000000010100000000100111" OR uut_a_5_4 /= "111100010111011000110010100" OR uut_a_5_5 /= "000110010010101100011110110" THEN
              FAIL <= '1';
              FAIL_NUM <= "01001110";
              state <= "11111101";
            ELSE
              state <= "01011100";
            END IF;
            uut_rst <= '0';
          WHEN "01011100" =>
            uut_coord_shift <= "1001";
            uut_x <= "110100011011";
            uut_y <= "110110111111";
            uut_fx <= "1010111011";
            uut_fy <= "1000101011";
            uut_ft <= "1001101110";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000110010110001" OR uut_a_0_1 /= "000000000110110101110110101" OR uut_a_0_2 /= "000000010110110110101011110" OR uut_a_0_3 /= "000000000000110010001101011" OR uut_a_0_4 /= "000000110110001000011010111" OR uut_a_0_5 /= "000010110100110101001010111" OR uut_a_1_0 /= "000000000000000001101101011" OR uut_a_1_1 /= "000000000001110110000000111" OR uut_a_1_2 /= "000000000110001010001111010" OR uut_a_1_3 /= "000000000000001101100010000" OR uut_a_1_4 /= "000000001110100101110001001" OR uut_a_1_5 /= "000000110000101111010101001" OR uut_a_2_0 /= "000000000000000101101101101" OR uut_a_2_1 /= "000000000110001010001111010" OR uut_a_2_2 /= "000000010100100100111111001" OR uut_a_2_3 /= "000000000000101101001101010" OR uut_a_2_4 /= "000000110000101111010101001" OR uut_a_2_5 /= "000010100010110100010111111" OR uut_a_3_0 /= "000000000000110010001101011" OR uut_a_3_1 /= "000000110110001000011010111" OR uut_a_3_2 /= "000010110100110101001010111" OR uut_a_3_3 /= "000000000110001101010001001" OR uut_a_3_4 /= "000110101100010011011101101" OR uut_a_3_5 /= "010110010110110010001011010" OR uut_a_4_0 /= "000000000000001101100010000" OR uut_a_4_1 /= "000000001110100101110001001" OR uut_a_4_2 /= "000000110000101111010101001" OR uut_a_4_3 /= "000000000001101011000100110" OR uut_a_4_4 /= "000001110011011100001111101" OR uut_a_4_5 /= "000110000001101001000001100" OR uut_a_5_0 /= "000000000000101101001101010" OR uut_a_5_1 /= "000000110000101111010101001" OR uut_a_5_2 /= "000010100010110100010111111" OR uut_a_5_3 /= "000000000101100101101100100" OR uut_a_5_4 /= "000110000001101001000001100" OR uut_a_5_5 /= "010100001000010000111011011" THEN
              FAIL <= '1';
              FAIL_NUM <= "01001111";
              state <= "11111101";
            ELSE
              state <= "01011101";
            END IF;
            uut_rst <= '0';
          WHEN "01011101" =>
            uut_coord_shift <= "1001";
            uut_x <= "000011101110";
            uut_y <= "001110000100";
            uut_fx <= "1101101011";
            uut_fy <= "1110100100";
            uut_ft <= "0111110000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000011111101000000100" OR uut_a_0_1 /= "001000010001101111001011011" OR uut_a_0_2 /= "110110110110111010101100110" OR uut_a_0_3 /= "111111111101110011110100111" OR uut_a_0_4 /= "111011011010100000101101010" OR uut_a_0_5 /= "000101000100001001101110100" OR uut_a_1_0 /= "000000000001000010001101111" OR uut_a_1_1 /= "000010001010101001000110001" OR uut_a_1_2 /= "111101100110110111110111001" OR uut_a_1_3 /= "111111111111011011010100000" OR uut_a_1_4 /= "111110110011001100000011110" OR uut_a_1_5 /= "000001010100110101100010111" OR uut_a_2_0 /= "111111111110110110110111010" OR uut_a_2_1 /= "111101100110110111110111001" OR uut_a_2_2 /= "000010101001001000000010000" OR uut_a_2_3 /= "000000000000101000100001001" OR uut_a_2_4 /= "000001010100110101100010111" OR uut_a_2_5 /= "111110100010010011001100000" OR uut_a_3_0 /= "111111111101110011110100111" OR uut_a_3_1 /= "111011011010100000101101010" OR uut_a_3_2 /= "000101000100001001101110100" OR uut_a_3_3 /= "000000000001001101101010010" OR uut_a_3_4 /= "000010100010100110011101100" OR uut_a_3_5 /= "111101001100011010010011000" OR uut_a_4_0 /= "111111111111011011010100000" OR uut_a_4_1 /= "111110110011001100000011110" OR uut_a_4_2 /= "000001010100110101100010111" OR uut_a_4_3 /= "000000000000010100010100110" OR uut_a_4_4 /= "000000101010100011100100001" OR uut_a_4_5 /= "111111010000111111111000011" OR uut_a_5_0 /= "000000000000101000100001001" OR uut_a_5_1 /= "000001010100110101100010111" OR uut_a_5_2 /= "111110100010010011001100000" OR uut_a_5_3 /= "111111111111101001100011010" OR uut_a_5_4 /= "111111010000111111111000011" OR uut_a_5_5 /= "000000110011111010011001100" THEN
              FAIL <= '1';
              FAIL_NUM <= "01010000";
              state <= "11111101";
            ELSE
              state <= "01011110";
            END IF;
            uut_rst <= '0';
          WHEN "01011110" =>
            uut_coord_shift <= "1001";
            uut_x <= "001110010000";
            uut_y <= "000101101001";
            uut_fx <= "0111110100";
            uut_fy <= "0100010001";
            uut_ft <= "1101011001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000010000010110100010" OR uut_a_0_1 /= "000011011011101110110000111" OR uut_a_0_2 /= "111100010100111100000111010" OR uut_a_0_3 /= "000000000010101101101101010" OR uut_a_0_4 /= "000100100011110001100000011" OR uut_a_0_5 /= "111011000111110111101100010" OR uut_a_1_0 /= "000000000000011011011101110" OR uut_a_1_1 /= "000000101110001000101000011" OR uut_a_1_2 /= "111111001110101001010111110" OR uut_a_1_3 /= "000000000000100100011110001" OR uut_a_1_4 /= "000000111101010000101101001" OR uut_a_1_5 /= "111110111110011101110000010" OR uut_a_2_0 /= "111111111111100010100111100" OR uut_a_2_1 /= "111111001110101001010111110" OR uut_a_2_2 /= "000000110100110010111111110" OR uut_a_2_3 /= "111111111111011000111110111" OR uut_a_2_4 /= "111110111110011101110000010" OR uut_a_2_5 /= "000001000110000110110111011" OR uut_a_3_0 /= "000000000010101101101101010" OR uut_a_3_1 /= "000100100011110001100000011" OR uut_a_3_2 /= "111011000111110111101100010" OR uut_a_3_3 /= "000000000011100110101010010" OR uut_a_3_4 /= "000110000011011011111101111" OR uut_a_3_5 /= "111001100001100010000101010" OR uut_a_4_0 /= "000000000000100100011110001" OR uut_a_4_1 /= "000000111101010000101101001" OR uut_a_4_2 /= "111110111110011101110000010" OR uut_a_4_3 /= "000000000000110000011011011" OR uut_a_4_4 /= "000001010001010110001011110" OR uut_a_4_5 /= "111110101000111110100101111" OR uut_a_5_0 /= "111111111111011000111110111" OR uut_a_5_1 /= "111110111110011101110000010" OR uut_a_5_2 /= "000001000110000110110111011" OR uut_a_5_3 /= "111111111111001100001100010" OR uut_a_5_4 /= "111110101000111110100101111" OR uut_a_5_5 /= "000001011101000101111110000" THEN
              FAIL <= '1';
              FAIL_NUM <= "01010001";
              state <= "11111101";
            ELSE
              state <= "01011111";
            END IF;
            uut_rst <= '0';
          WHEN "01011111" =>
            uut_coord_shift <= "1001";
            uut_x <= "000101001100";
            uut_y <= "110111110101";
            uut_fx <= "1100101111";
            uut_fy <= "0010111001";
            uut_ft <= "0000011101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000010001010001100" OR uut_a_0_1 /= "111110101000110100010111010" OR uut_a_0_2 /= "000000111110010110011000111" OR uut_a_0_3 /= "111111111111010010100010101" OR uut_a_0_4 /= "000011100101011011010000001" OR uut_a_0_5 /= "111101011011111010111110011" OR uut_a_1_0 /= "111111111111110101000110100" OR uut_a_1_1 /= "000000110110111111111101110" OR uut_a_1_2 /= "111111011000101010101000000" OR uut_a_1_3 /= "000000000000011100101011011" OR uut_a_1_4 /= "111101101111010000111011101" OR uut_a_1_5 /= "000001100111100000101010111" OR uut_a_2_0 /= "000000000000000111110010110" OR uut_a_2_1 /= "111111011000101010101000000" OR uut_a_2_2 /= "000000011100001000010110100" OR uut_a_2_3 /= "111111111111101011011111010" OR uut_a_2_4 /= "000001100111100000101010111" OR uut_a_2_5 /= "111110110101111110001110111" OR uut_a_3_0 /= "111111111111010010100010101" OR uut_a_3_1 /= "000011100101011011010000001" OR uut_a_3_2 /= "111101011011111010111110011" OR uut_a_3_3 /= "000000000001110111101000010" OR uut_a_3_4 /= "110110100100001111110111010" OR uut_a_3_5 /= "000110101111110010010001110" OR uut_a_4_0 /= "000000000000011100101011011" OR uut_a_4_1 /= "111101101111010000111011101" OR uut_a_4_2 /= "000001100111100000101010111" OR uut_a_4_3 /= "111111111110110100100001111" OR uut_a_4_4 /= "000101111100111000011111100" OR uut_a_4_5 /= "111011101111100110101010000" OR uut_a_5_0 /= "111111111111101011011111010" OR uut_a_5_1 /= "000001100111100000101010111" OR uut_a_5_2 /= "111110110101111110001110111" OR uut_a_5_3 /= "000000000000110101111110010" OR uut_a_5_4 /= "111011101111100110101010000" OR uut_a_5_5 /= "000011000010110011110011110" THEN
              FAIL <= '1';
              FAIL_NUM <= "01010010";
              state <= "11111101";
            ELSE
              state <= "01100000";
            END IF;
            uut_rst <= '0';
          WHEN "01100000" =>
            uut_coord_shift <= "1001";
            uut_x <= "111101001011";
            uut_y <= "000011010010";
            uut_fx <= "0100000001";
            uut_fy <= "0001010110";
            uut_ft <= "0000110101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000011010101111001000" OR uut_a_0_1 /= "000011110010010011000100100" OR uut_a_0_2 /= "101110101111011101001001100" OR uut_a_0_3 /= "111111111110010010010100000" OR uut_a_0_4 /= "111110000011101111101010000" OR uut_a_0_5 /= "001000110110011011101110000" OR uut_a_1_0 /= "000000000000011110010010011" OR uut_a_1_1 /= "000000100010010011110100110" OR uut_a_1_2 /= "111101100011100110000100001" OR uut_a_1_3 /= "111111111111110000011101111" OR uut_a_1_4 /= "111111101110011001111011111" OR uut_a_1_5 /= "000001010000001101010011001" OR uut_a_2_0 /= "111111111101110101111011101" OR uut_a_2_1 /= "111101100011100110000100001" OR uut_a_2_2 /= "001011001000111111011111110" OR uut_a_2_3 /= "000000000001000110110011011" OR uut_a_2_4 /= "000001010000001101010011001" OR uut_a_2_5 /= "111010010010010111001110110" OR uut_a_3_0 /= "111111111110010010010100000" OR uut_a_3_1 /= "111110000011101111101010000" OR uut_a_3_2 /= "001000110110011011101110000" OR uut_a_3_3 /= "000000000000111000010000000" OR uut_a_3_4 /= "000000111111101110001000000" OR uut_a_3_5 /= "111011011101100001011000000" OR uut_a_4_0 /= "111111111111110000011101111" OR uut_a_4_1 /= "111111101110011001111011111" OR uut_a_4_2 /= "000001010000001101010011001" OR uut_a_4_3 /= "000000000000000111111101110" OR uut_a_4_4 /= "000000001001000001011110000" OR uut_a_4_5 /= "111111010110110111100010011" OR uut_a_5_0 /= "000000000001000110110011011" OR uut_a_5_1 /= "000001010000001101010011001" OR uut_a_5_2 /= "111010010010010111001110110" OR uut_a_5_3 /= "111111111111011011101100001" OR uut_a_5_4 /= "111111010110110111100010011" OR uut_a_5_5 /= "000010111011100000011001001" THEN
              FAIL <= '1';
              FAIL_NUM <= "01010011";
              state <= "11111101";
            ELSE
              state <= "01100001";
            END IF;
            uut_rst <= '0';
          WHEN "01100001" =>
            uut_coord_shift <= "1001";
            uut_x <= "000010101011";
            uut_y <= "000000011000";
            uut_fx <= "1001010101";
            uut_fy <= "0011100001";
            uut_ft <= "0111111100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000010101101111010010" OR uut_a_0_1 /= "110100000000010110011000011" OR uut_a_0_2 /= "111010100001011101100101110" OR uut_a_0_3 /= "111111111111000101000100011" OR uut_a_0_4 /= "000100000100001000001100000" OR uut_a_0_5 /= "000001110110110010001011101" OR uut_a_1_0 /= "111111111110100000000010110" OR uut_a_1_1 /= "000110100111100011101001101" OR uut_a_1_2 /= "000011000001011010010111000" OR uut_a_1_3 /= "000000000000100000100001000" OR uut_a_1_4 /= "111101110000011110001110110" OR uut_a_1_5 /= "111110111110011101011011111" OR uut_a_2_0 /= "111111111111010100001011101" OR uut_a_2_1 /= "000011000001011010010111000" OR uut_a_2_2 /= "000001011000010100011010110" OR uut_a_2_3 /= "000000000000001110110110010" OR uut_a_2_4 /= "111110111110011101011011111" OR uut_a_2_5 /= "111111100010000100100110110" OR uut_a_3_0 /= "111111111111000101000100011" OR uut_a_3_1 /= "000100000100001000001100000" OR uut_a_3_2 /= "000001110110110010001011101" OR uut_a_3_3 /= "000000000000010011111110000" OR uut_a_3_4 /= "111110100111110110100011010" OR uut_a_3_5 /= "111111010111101111111001111" OR uut_a_4_0 /= "000000000000100000100001000" OR uut_a_4_1 /= "111101110000011110001110110" OR uut_a_4_2 /= "111110111110011101011011111" OR uut_a_4_3 /= "111111111111110100111110110" OR uut_a_4_4 /= "000000110000101000101101100" OR uut_a_4_5 /= "000000010110001101011000010" OR uut_a_5_0 /= "000000000000001110110110010" OR uut_a_5_1 /= "111110111110011101011011111" OR uut_a_5_2 /= "111111100010000100100110110" OR uut_a_5_3 /= "111111111111111010111101111" OR uut_a_5_4 /= "000000010110001101011000010" OR uut_a_5_5 /= "000000001010001001000011100" THEN
              FAIL <= '1';
              FAIL_NUM <= "01010100";
              state <= "11111101";
            ELSE
              state <= "01100010";
            END IF;
            uut_rst <= '0';
          WHEN "01100010" =>
            uut_coord_shift <= "1001";
            uut_x <= "111011010111";
            uut_y <= "001111000101";
            uut_fx <= "1101100011";
            uut_fy <= "0110001100";
            uut_ft <= "1111010010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000010111110001000" OR uut_a_0_1 /= "111101010011001001000110100" OR uut_a_0_2 /= "000001010100110110011100100" OR uut_a_0_3 /= "111111111111100111000001000" OR uut_a_0_4 /= "000010110101101110001110100" OR uut_a_0_5 /= "111110100110110011000100100" OR uut_a_1_0 /= "111111111111101010011001001" OR uut_a_1_1 /= "000010011101001010001010011" OR uut_a_1_2 /= "111110110010110110101111111" OR uut_a_1_3 /= "000000000000010110101101110" OR uut_a_1_4 /= "111101011010110010000010001" OR uut_a_1_5 /= "000001010001000110011100010" OR uut_a_2_0 /= "000000000000001010100110110" OR uut_a_2_1 /= "111110110010110110101111111" OR uut_a_2_2 /= "000000100101110111100011000" OR uut_a_2_3 /= "111111111111110100110110011" OR uut_a_2_4 /= "000001010001000110011100010" OR uut_a_2_5 /= "111111011000001100001010101" OR uut_a_3_0 /= "111111111111100111000001000" OR uut_a_3_1 /= "000010110101101110001110100" OR uut_a_3_2 /= "111110100110110011000100100" OR uut_a_3_3 /= "000000000000011010010001000" OR uut_a_3_4 /= "111101000000111101010110100" OR uut_a_3_5 /= "000001011101110001101100100" OR uut_a_4_0 /= "000000000000010110101101110" OR uut_a_4_1 /= "111101011010110010000010001" OR uut_a_4_2 /= "000001010001000110011100010" OR uut_a_4_3 /= "111111111111101000000111101" OR uut_a_4_4 /= "000010101101101100001110000" OR uut_a_4_5 /= "111110101010101111011000010" OR uut_a_5_0 /= "111111111111110100110110011" OR uut_a_5_1 /= "000001010001000110011100010" OR uut_a_5_2 /= "111111011000001100001010101" OR uut_a_5_3 /= "000000000000001011101110001" OR uut_a_5_4 /= "111110101010101111011000010" OR uut_a_5_5 /= "000000101001110110011111011" THEN
              FAIL <= '1';
              FAIL_NUM <= "01010101";
              state <= "11111101";
            ELSE
              state <= "01100011";
            END IF;
            uut_rst <= '0';
          WHEN "01100011" =>
            uut_coord_shift <= "1001";
            uut_x <= "111101001111";
            uut_y <= "110110111110";
            uut_fx <= "1010000001";
            uut_fy <= "1100111100";
            uut_ft <= "0011101000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000010101100010001000" OR uut_a_0_1 /= "000101011101111010100010000" OR uut_a_0_2 /= "101011011010011011111110100" OR uut_a_0_3 /= "000000000001111110010101000" OR uut_a_0_4 /= "000100000000100110101010000" OR uut_a_0_5 /= "110000111001110010011000100" OR uut_a_1_0 /= "000000000000101011101111010" OR uut_a_1_1 /= "000001011000110110000111001" OR uut_a_1_2 /= "111010110001011101100110100" OR uut_a_1_3 /= "000000000000100000000100110" OR uut_a_1_4 /= "000001000001001001110100001" OR uut_a_1_5 /= "111100001010101011000010101" OR uut_a_2_0 /= "111111111101011011010011011" OR uut_a_2_1 /= "111010110001011101100110100" OR uut_a_2_2 /= "010011101011101010011000001" OR uut_a_2_3 /= "111111111110000111001110010" OR uut_a_2_4 /= "111100001010101011000010101" OR uut_a_2_5 /= "001110011011110000001001001" OR uut_a_3_0 /= "000000000001111110010101000" OR uut_a_3_1 /= "000100000000100110101010000" OR uut_a_3_2 /= "110000111001110010011000100" OR uut_a_3_3 /= "000000000001011100101001000" OR uut_a_3_4 /= "000010111100001011010010000" OR uut_a_3_5 /= "110100111011011100011010100" OR uut_a_4_0 /= "000000000000100000000100110" OR uut_a_4_1 /= "000001000001001001110100001" OR uut_a_4_2 /= "111100001010101011000010101" OR uut_a_4_3 /= "000000000000010111100001011" OR uut_a_4_4 /= "000000101111110001110111010" OR uut_a_4_5 /= "111101001100000101111101101" OR uut_a_5_0 /= "111111111110000111001110010" OR uut_a_5_1 /= "111100001010101011000010101" OR uut_a_5_2 /= "001110011011110000001001001" OR uut_a_5_3 /= "111111111110100111011011100" OR uut_a_5_4 /= "111101001100000101111101101" OR uut_a_5_5 /= "001010100101011010110001011" THEN
              FAIL <= '1';
              FAIL_NUM <= "01010110";
              state <= "11111101";
            ELSE
              state <= "01100100";
            END IF;
            uut_rst <= '0';
          WHEN "01100100" =>
            uut_coord_shift <= "1010";
            uut_x <= "010010000110";
            uut_y <= "001100011001";
            uut_fx <= "1000001010";
            uut_fy <= "0101011111";
            uut_ft <= "0110110000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000001110000100000" OR uut_a_0_1 /= "000001000110011011000010000" OR uut_a_0_2 /= "111111100101110110100100000" OR uut_a_0_3 /= "000000000000001001000001100" OR uut_a_0_4 /= "000000101101001100000000110" OR uut_a_0_5 /= "111111101111001110001101100" OR uut_a_1_0 /= "000000000000001000110011011" OR uut_a_1_1 /= "000000101100000101010010111" OR uut_a_1_2 /= "111111101111101000011101111" OR uut_a_1_3 /= "000000000000000101101001100" OR uut_a_1_4 /= "000000011100010010010101001" OR uut_a_1_5 /= "111111110101011111110101010" OR uut_a_2_0 /= "111111111111111100101110110" OR uut_a_2_1 /= "111111101111101000011101111" OR uut_a_2_2 /= "000000000110000100111100011" OR uut_a_2_3 /= "111111111111111101111001110" OR uut_a_2_4 /= "111111110101011111110101010" OR uut_a_2_5 /= "000000000011111001100100100" OR uut_a_3_0 /= "000000000000001001000001100" OR uut_a_3_1 /= "000000101101001100000000110" OR uut_a_3_2 /= "111111101111001110001101100" OR uut_a_3_3 /= "000000000000000101110010100" OR uut_a_3_4 /= "000000011100111111101101010" OR uut_a_3_5 /= "111111110101001110111111000" OR uut_a_4_0 /= "000000000000000101101001100" OR uut_a_4_1 /= "000000011100010010010101001" OR uut_a_4_2 /= "111111110101011111110101010" OR uut_a_4_3 /= "000000000000000011100111111" OR uut_a_4_4 /= "000000010010001001101000010" OR uut_a_4_5 /= "111111111001010000101100010" OR uut_a_5_0 /= "111111111111111101111001110" OR uut_a_5_1 /= "111111110101011111110101010" OR uut_a_5_2 /= "000000000011111001100100100" OR uut_a_5_3 /= "111111111111111110101001110" OR uut_a_5_4 /= "111111111001010000101100010" OR uut_a_5_5 /= "000000000010100000001001000" THEN
              FAIL <= '1';
              FAIL_NUM <= "01010111";
              state <= "11111101";
            ELSE
              state <= "01100101";
            END IF;
            uut_rst <= '0';
          WHEN "01100101" =>
            uut_coord_shift <= "1010";
            uut_x <= "010001010101";
            uut_y <= "100010101111";
            uut_fx <= "1110000011";
            uut_fy <= "0011010001";
            uut_ft <= "0011101011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000010011100010" OR uut_a_0_1 /= "111111110111001110011110100" OR uut_a_0_2 /= "111111110110001100100011110" OR uut_a_0_3 /= "000000000000001101100111111" OR uut_a_0_4 /= "111111001111000010101100110" OR uut_a_0_5 /= "111111001001010010111000001" OR uut_a_1_0 /= "111111111111111110111001110" OR uut_a_1_1 /= "000000000011111100001111110" OR uut_a_1_2 /= "000000000100011001110110111" OR uut_a_1_3 /= "111111111111111001111000010" OR uut_a_1_4 /= "000000010101111111100010011" OR uut_a_1_5 /= "000000011000100100110001010" OR uut_a_2_0 /= "111111111111111110110001100" OR uut_a_2_1 /= "000000000100011001110110111" OR uut_a_2_2 /= "000000000100111010111100100" OR uut_a_2_3 /= "111111111111111001001010010" OR uut_a_2_4 /= "000000011000100100110001010" OR uut_a_2_5 /= "000000011011011101011001100" OR uut_a_3_0 /= "000000000000001101100111111" OR uut_a_3_1 /= "111111001111000010101100110" OR uut_a_3_2 /= "111111001001010010111000001" OR uut_a_3_3 /= "000000000001001100000001000" OR uut_a_3_4 /= "111011101110110100001011101" OR uut_a_3_5 /= "111011001110101111101110111" OR uut_a_4_0 /= "111111111111111001111000010" OR uut_a_4_1 /= "000000010101111111100010011" OR uut_a_4_2 /= "000000011000100100110001010" OR uut_a_4_3 /= "111111111111011101110110100" OR uut_a_4_4 /= "000001111010101110000011110" OR uut_a_4_5 /= "000010001001001000000011101" OR uut_a_5_0 /= "111111111111111001001010010" OR uut_a_5_1 /= "000000011000100100110001010" OR uut_a_5_2 /= "000000011011011101011001100" OR uut_a_5_3 /= "111111111111011001110101111" OR uut_a_5_4 /= "000010001001001000000011101" OR uut_a_5_5 /= "000010011001001110010010100" THEN
              FAIL <= '1';
              FAIL_NUM <= "01011000";
              state <= "11111101";
            ELSE
              state <= "01100110";
            END IF;
            uut_rst <= '0';
          WHEN "01100110" =>
            uut_coord_shift <= "1010";
            uut_x <= "101110010111";
            uut_y <= "110001001111";
            uut_fx <= "0010110001";
            uut_fy <= "1111101001";
            uut_ft <= "0001111111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000001010101100" OR uut_a_0_1 /= "000000001010011001000111010" OR uut_a_0_2 /= "111111110101111100111100011" OR uut_a_0_3 /= "111111111111110000101101110" OR uut_a_0_4 /= "111110001001001100000111101" OR uut_a_0_5 /= "000001110010110111101100001" OR uut_a_1_0 /= "000000000000000001010011001" OR uut_a_1_1 /= "000000001010000110010001110" OR uut_a_1_2 /= "111111110110001111001001111" OR uut_a_1_3 /= "111111111111110001001001100" OR uut_a_1_4 /= "111110001100100011011101110" OR uut_a_1_5 /= "000001101111100111011111001" OR uut_a_2_0 /= "111111111111111110101111100" OR uut_a_2_1 /= "111111110110001111001001111" OR uut_a_2_2 /= "000000001001011100000111101" OR uut_a_2_3 /= "000000000000001110010110111" OR uut_a_2_4 /= "000001101111100111011111001" OR uut_a_2_5 /= "111110010100000101011011100" OR uut_a_3_0 /= "111111111111110000101101110" OR uut_a_3_1 /= "111110001001001100000111101" OR uut_a_3_2 /= "000001110010110111101100001" OR uut_a_3_3 /= "000000000010101110101111000" OR uut_a_3_4 /= "010101001110010010110101100" OR uut_a_3_5 /= "101011011110110000010010111" OR uut_a_4_0 /= "111111111111110001001001100" OR uut_a_4_1 /= "111110001100100011011101110" OR uut_a_4_2 /= "000001101111100111011111001" OR uut_a_4_3 /= "000000000010101001110010010" OR uut_a_4_4 /= "010100100111110100111011011" OR uut_a_4_5 /= "101100000011111100100011011" OR uut_a_5_0 /= "000000000000001110010110111" OR uut_a_5_1 /= "000001101111100111011111001" OR uut_a_5_2 /= "111110010100000101011011100" OR uut_a_5_3 /= "111111111101011011110110000" OR uut_a_5_4 /= "101100000011111100100011011" OR uut_a_5_5 /= "010011010001101110111000001" THEN
              FAIL <= '1';
              FAIL_NUM <= "01011001";
              state <= "11111101";
            ELSE
              state <= "01100111";
            END IF;
            uut_rst <= '0';
          WHEN "01100111" =>
            uut_coord_shift <= "1010";
            uut_x <= "101111001001";
            uut_y <= "101011010110";
            uut_fx <= "0101010010";
            uut_fy <= "0100010001";
            uut_ft <= "0110111101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000011000101110000010" OR uut_a_0_1 /= "011000001010011111110101001" OR uut_a_0_2 /= "101010100111001011000001010" OR uut_a_0_3 /= "111111111100100111010110011" OR uut_a_0_4 /= "100101100001101110011110101" OR uut_a_0_5 /= "010111011011101000000111111" OR uut_a_1_0 /= "000000000011000001010011111" OR uut_a_1_1 /= "010111100111110000101111010" OR uut_a_1_2 /= "101011000101111010101101011" OR uut_a_1_3 /= "111111111100101100001101110" OR uut_a_1_4 /= "100110000111110001111111110" OR uut_a_1_5 /= "010110111001111100011010001" OR uut_a_2_0 /= "111111111101010100111001011" OR uut_a_2_1 /= "101011000101111010101101011" OR uut_a_2_2 /= "010010100000010110110101110" OR uut_a_2_3 /= "000000000010111011011101000" OR uut_a_2_4 /= "010110111001111100011010001" OR uut_a_2_5 /= "101011101110011110001010001" OR uut_a_3_0 /= "111111111100100111010110011" OR uut_a_3_1 /= "100101100001101110011110101" OR uut_a_3_2 /= "010111011011101000000111111" OR uut_a_3_3 /= "000000000011101101010110100" OR uut_a_3_4 /= "011101000000001010111100100" OR uut_a_3_5 /= "100110010101000100110100110" OR uut_a_4_0 /= "111111111100101100001101110" OR uut_a_4_1 /= "100110000111110001111111110" OR uut_a_4_2 /= "010110111001111100011010001" OR uut_a_4_3 /= "000000000011101000000001010" OR uut_a_4_4 /= "011100010110011110101100110" OR uut_a_4_5 /= "100110111001111110100001111" OR uut_a_5_0 /= "000000000010111011011101000" OR uut_a_5_1 /= "010110111001111100011010001" OR uut_a_5_2 /= "101011101110011110001010001" OR uut_a_5_3 /= "111111111100110010101000100" OR uut_a_5_4 /= "100110111001111110100001111" OR uut_a_5_5 /= "010110001101100000111100110" THEN
              FAIL <= '1';
              FAIL_NUM <= "01011010";
              state <= "11111101";
            ELSE
              state <= "01101000";
            END IF;
            uut_rst <= '0';
          WHEN "01101000" =>
            uut_coord_shift <= "1010";
            uut_x <= "100110111010";
            uut_y <= "101011101011";
            uut_fx <= "1001100101";
            uut_fy <= "1111110110";
            uut_ft <= "1011000110";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000010011000010111100" OR uut_a_0_1 /= "001010110011100110111100111" OR uut_a_0_2 /= "000001010010001000101100111" OR uut_a_0_3 /= "000000000010011101110001001" OR uut_a_0_4 /= "001011001100000111110000111" OR uut_a_0_5 /= "000001010101000011000000111" OR uut_a_1_0 /= "000000000001010110011100110" OR uut_a_1_1 /= "000110001000011010000010011" OR uut_a_1_2 /= "000000101110100110100011111" OR uut_a_1_3 /= "000000000001011001100000111" OR uut_a_1_4 /= "000110010110010100001001111" OR uut_a_1_5 /= "000000110000010000010001011" OR uut_a_2_0 /= "000000000000001010010001000" OR uut_a_2_1 /= "000000101110100110100011111" OR uut_a_2_2 /= "000000000101100010001101100" OR uut_a_2_3 /= "000000000000001010101000011" OR uut_a_2_4 /= "000000110000010000010001011" OR uut_a_2_5 /= "000000000101101110110001000" OR uut_a_3_0 /= "000000000010011101110001001" OR uut_a_3_1 /= "001011001100000111110000111" OR uut_a_3_2 /= "000001010101000011000000111" OR uut_a_3_3 /= "000000000010100011010111000" OR uut_a_3_4 /= "001011100101100000001011101" OR uut_a_3_5 /= "000001011000000011111011101" OR uut_a_4_0 /= "000000000001011001100000111" OR uut_a_4_1 /= "000110010110010100001001111" OR uut_a_4_2 /= "000000110000010000010001011" OR uut_a_4_3 /= "000000000001011100101100000" OR uut_a_4_4 /= "000110100100101101110100100" OR uut_a_4_5 /= "000000110001111101101110110" OR uut_a_5_0 /= "000000000000001010101000011" OR uut_a_5_1 /= "000000110000010000010001011" OR uut_a_5_2 /= "000000000101101110110001000" OR uut_a_5_3 /= "000000000000001011000000011" OR uut_a_5_4 /= "000000110001111101101110110" OR uut_a_5_5 /= "000000000101111011110000111" THEN
              FAIL <= '1';
              FAIL_NUM <= "01011011";
              state <= "11111101";
            ELSE
              state <= "01101001";
            END IF;
            uut_rst <= '0';
          WHEN "01101001" =>
            uut_coord_shift <= "1010";
            uut_x <= "011001010101";
            uut_y <= "100110010110";
            uut_fx <= "1000101101";
            uut_fy <= "0000111011";
            uut_ft <= "0100010111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001100111001001100" OR uut_a_0_1 /= "110110101010110111001001000" OR uut_a_0_2 /= "111000101111000001011001001" OR uut_a_0_3 /= "000000000010010100110110100" OR uut_a_0_4 /= "110010100010010010001000100" OR uut_a_0_5 /= "110101100001000000000010101" OR uut_a_1_0 /= "111111111110110101010110111" OR uut_a_1_1 /= "000110110000000110111110001" OR uut_a_1_2 /= "000101010000011110010011011" OR uut_a_1_3 /= "111111111110010100010010010" OR uut_a_1_4 /= "001001101111100100010000001" OR uut_a_1_5 /= "000111100101100011101010000" OR uut_a_2_0 /= "111111111111000101111000001" OR uut_a_2_1 /= "000101010000011110010011011" OR uut_a_2_2 /= "000100000110000000010001101" OR uut_a_2_3 /= "111111111110101100001000000" OR uut_a_2_4 /= "000111100101100011101010000" OR uut_a_2_5 /= "000101111010000101111010011" OR uut_a_3_0 /= "000000000010010100110110100" OR uut_a_3_1 /= "110010100010010010001000100" OR uut_a_3_2 /= "110101100001000000000010101" OR uut_a_3_3 /= "000000000011010110110011100" OR uut_a_3_4 /= "101100100100011110100000000" OR uut_a_3_5 /= "110000110111101100100100001" OR uut_a_4_0 /= "111111111110010100010010010" OR uut_a_4_1 /= "001001101111100100010000001" OR uut_a_4_2 /= "000111100101100011101010000" OR uut_a_4_3 /= "111111111101100100100011110" OR uut_a_4_4 /= "001110000011110110101011011" OR uut_a_4_5 /= "001010111100101100100100000" OR uut_a_5_0 /= "111111111110101100001000000" OR uut_a_5_1 /= "000111100101100011101010000" OR uut_a_5_2 /= "000101111010000101111010011" OR uut_a_5_3 /= "111111111110000110111101100" OR uut_a_5_4 /= "001010111100101100100100000" OR uut_a_5_5 /= "001000100001100111011100110" THEN
              FAIL <= '1';
              FAIL_NUM <= "01011100";
              state <= "11111101";
            ELSE
              state <= "01101010";
            END IF;
            uut_rst <= '0';
          WHEN "01101010" =>
            uut_coord_shift <= "1010";
            uut_x <= "110011111110";
            uut_y <= "101011011110";
            uut_fx <= "1101011011";
            uut_fy <= "1011010111";
            uut_ft <= "0000001010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000010101101011100" OR uut_a_0_1 /= "000000101000010011111111111" OR uut_a_0_2 /= "000010011000011100010011001" OR uut_a_0_3 /= "000000000000001101011000110" OR uut_a_0_4 /= "000000011000111001000001010" OR uut_a_0_5 /= "000001011110001000000001100" OR uut_a_1_0 /= "000000000000000101000010011" OR uut_a_1_1 /= "000000001001010111101001011" OR uut_a_1_2 /= "000000100011011011100100111" OR uut_a_1_3 /= "000000000000000011000111001" OR uut_a_1_4 /= "000000000101110010010000001" OR uut_a_1_5 /= "000000010101111000000111010" OR uut_a_2_0 /= "000000000000010011000011100" OR uut_a_2_1 /= "000000100011011011100100111" OR uut_a_2_2 /= "000010000101111110110111110" OR uut_a_2_3 /= "000000000000001011110001000" OR uut_a_2_4 /= "000000010101111000000111010" OR uut_a_2_5 /= "000001010010101110100011010" OR uut_a_3_0 /= "000000000000001101011000110" OR uut_a_3_1 /= "000000011000111001000001010" OR uut_a_3_2 /= "000001011110001000000001100" OR uut_a_3_3 /= "000000000000001000010001000" OR uut_a_3_4 /= "000000001111010111100111000" OR uut_a_3_5 /= "000000111010000111100010000" OR uut_a_4_0 /= "000000000000000011000111001" OR uut_a_4_1 /= "000000000101110010010000001" OR uut_a_4_2 /= "000000010101111000000111010" OR uut_a_4_3 /= "000000000000000001111010111" OR uut_a_4_4 /= "000000000011100100100111001" OR uut_a_4_5 /= "000000001101100000100000000" OR uut_a_5_0 /= "000000000000001011110001000" OR uut_a_5_1 /= "000000010101111000000111010" OR uut_a_5_2 /= "000001010010101110100011010" OR uut_a_5_3 /= "000000000000000111010000111" OR uut_a_5_4 /= "000000001101100000100000000" OR uut_a_5_5 /= "000000110011000101000111101" THEN
              FAIL <= '1';
              FAIL_NUM <= "01011101";
              state <= "11111101";
            ELSE
              state <= "01101011";
            END IF;
            uut_rst <= '0';
          WHEN "01101011" =>
            uut_coord_shift <= "1010";
            uut_x <= "011010000000";
            uut_y <= "001000010000";
            uut_fx <= "1001101000";
            uut_fy <= "1110010000";
            uut_ft <= "1000111000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000011110100001001000" OR uut_a_0_1 /= "011011001011100000001000000" OR uut_a_0_2 /= "001010110000100011011000100" OR uut_a_0_3 /= "000000000010000101010011010" OR uut_a_0_4 /= "001110110101110001001010000" OR uut_a_0_5 /= "000101110111111100110010101" OR uut_a_1_0 /= "000000000011011001011100000" OR uut_a_1_1 /= "011000001101001111100111001" OR uut_a_1_2 /= "001001100101001111100000110" OR uut_a_1_3 /= "000000000001110110101110001" OR uut_a_1_4 /= "001101001101111000110001111" OR uut_a_1_5 /= "000101001110110101001001000" OR uut_a_2_0 /= "000000000001010110000100011" OR uut_a_2_1 /= "001001100101001111100000110" OR uut_a_2_2 /= "000011110010101111011110010" OR uut_a_2_3 /= "000000000000101110111111100" OR uut_a_2_4 /= "000101001110110101001001000" OR uut_a_2_5 /= "000010000100100010010111100" OR uut_a_3_0 /= "000000000010000101010011010" OR uut_a_3_1 /= "001110110101110001001010000" OR uut_a_3_2 /= "000101110111111100110010101" OR uut_a_3_3 /= "000000000001001000110010000" OR uut_a_3_4 /= "001000000110100100101100100" OR uut_a_3_5 /= "000011001101010001001100010" OR uut_a_4_0 /= "000000000001110110101110001" OR uut_a_4_1 /= "001101001101111000110001111" OR uut_a_4_2 /= "000101001110110101001001000" OR uut_a_4_3 /= "000000000001000000110100100" OR uut_a_4_4 /= "000111001101110110101011101" OR uut_a_4_5 /= "000010110110110100010011111" OR uut_a_5_0 /= "000000000000101110111111100" OR uut_a_5_1 /= "000101001110110101001001000" OR uut_a_5_2 /= "000010000100100010010111100" OR uut_a_5_3 /= "000000000000011001101010001" OR uut_a_5_4 /= "000010110110110100010011111" OR uut_a_5_5 /= "000001001000010111010111111" THEN
              FAIL <= '1';
              FAIL_NUM <= "01011110";
              state <= "11111101";
            ELSE
              state <= "01101100";
            END IF;
            uut_rst <= '0';
          WHEN "01101100" =>
            uut_coord_shift <= "1010";
            uut_x <= "000000000101";
            uut_y <= "111011101001";
            uut_fx <= "0111111110";
            uut_fy <= "0100111111";
            uut_ft <= "1111110001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000101010101010000" OR uut_a_0_1 /= "000001101110101001000110011" OR uut_a_0_2 /= "111101010001101101001000101" OR uut_a_0_3 /= "111111111111011010001111011" OR uut_a_0_4 /= "111110011110000100000010101" OR uut_a_0_5 /= "000010011010010001111011000" OR uut_a_1_0 /= "000000000000001101110101001" OR uut_a_1_1 /= "000000100011110111110100110" OR uut_a_1_2 /= "111111000111011111011000100" OR uut_a_1_3 /= "111111111111110011110000100" OR uut_a_1_4 /= "111111100000001111110011110" OR uut_a_1_5 /= "000000110010000001010011111" OR uut_a_2_0 /= "111111111111101010001101101" OR uut_a_2_1 /= "111111000111011111011000100" OR uut_a_2_2 /= "000001011001000001010000101" OR uut_a_2_3 /= "000000000000010011010010001" OR uut_a_2_4 /= "000000110010000001010011111" OR uut_a_2_5 /= "111110110001001100111110001" OR uut_a_3_0 /= "111111111111011010001111011" OR uut_a_3_1 /= "111110011110000100000010101" OR uut_a_3_2 /= "000010011010010001111011000" OR uut_a_3_3 /= "000000000000100001011011000" OR uut_a_3_4 /= "000001010110101100001100011" OR uut_a_3_5 /= "111101110111011011111011001" OR uut_a_4_0 /= "111111111111110011110000100" OR uut_a_4_1 /= "111111100000001111110011110" OR uut_a_4_2 /= "000000110010000001010011111" OR uut_a_4_3 /= "000000000000001010110101100" OR uut_a_4_4 /= "000000011100000110110101000" OR uut_a_4_5 /= "111111010011101110010011011" OR uut_a_5_0 /= "000000000000010011010010001" OR uut_a_5_1 /= "000000110010000001010011111" OR uut_a_5_2 /= "111110110001001100111110001" OR uut_a_5_3 /= "111111111111101110111011011" OR uut_a_5_4 /= "111111010011101110010011011" OR uut_a_5_5 /= "000001000101101111111011001" THEN
              FAIL <= '1';
              FAIL_NUM <= "01011111";
              state <= "11111101";
            ELSE
              state <= "01101101";
            END IF;
            uut_rst <= '0';
          WHEN "01101101" =>
            uut_coord_shift <= "1010";
            uut_x <= "011001001111";
            uut_y <= "101000110100";
            uut_fx <= "1110001111";
            uut_fy <= "0110110110";
            uut_ft <= "0110101100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001000000100000000" OR uut_a_0_1 /= "111110100100110010101010010" OR uut_a_0_2 /= "000001101001110100100110100" OR uut_a_0_3 /= "000000000000010101100101011" OR uut_a_0_4 /= "111111100001011110101001100" OR uut_a_0_5 /= "000000100011011010010100011" OR uut_a_1_0 /= "111111111111110100100110010" OR uut_a_1_1 /= "000000010000000111110010111" OR uut_a_1_2 /= "111111101101010010111000111" OR uut_a_1_3 /= "111111111111111100001011110" OR uut_a_1_4 /= "000000000101011001010001010" OR uut_a_1_5 /= "111111111001101111011010010" OR uut_a_2_0 /= "000000000000001101001110100" OR uut_a_2_1 /= "111111101101010010111000111" OR uut_a_2_2 /= "000000010101101100111010011" OR uut_a_2_3 /= "000000000000000100011011010" OR uut_a_2_4 /= "111111111001101111011010010" OR uut_a_2_5 /= "000000000111010000110001011" OR uut_a_3_0 /= "000000000000010101100101011" OR uut_a_3_1 /= "111111100001011110101001100" OR uut_a_3_2 /= "000000100011011010010100011" OR uut_a_3_3 /= "000000000000000111001110010" OR uut_a_3_4 /= "111111110101110010010110011" OR uut_a_3_5 /= "000000001011110110011000010" OR uut_a_4_0 /= "111111111111111100001011110" OR uut_a_4_1 /= "000000000101011001010001010" OR uut_a_4_2 /= "111111111001101111011010010" OR uut_a_4_3 /= "111111111111111110101110010" OR uut_a_4_4 /= "000000000001110011100010011" OR uut_a_4_5 /= "111111111101111001111100110" OR uut_a_5_0 /= "000000000000000100011011010" OR uut_a_5_1 /= "111111111001101111011010010" OR uut_a_5_2 /= "000000000111010000110001011" OR uut_a_5_3 /= "000000000000000001011110110" OR uut_a_5_4 /= "111111111101111001111100110" OR uut_a_5_5 /= "000000000010011011100001101" THEN
              FAIL <= '1';
              FAIL_NUM <= "01100000";
              state <= "11111101";
            ELSE
              state <= "01101110";
            END IF;
            uut_rst <= '0';
          WHEN "01101110" =>
            uut_coord_shift <= "1010";
            uut_x <= "001101101010";
            uut_y <= "000111100100";
            uut_fx <= "1101100000";
            uut_fy <= "0110111110";
            uut_ft <= "1010000000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000010110010000011100" OR uut_a_0_1 /= "000011101101110111110000100" OR uut_a_0_2 /= "000000100001011000101010110" OR uut_a_0_3 /= "111111111110100010001011010" OR uut_a_0_4 /= "111110000010101010000111001" OR uut_a_0_5 /= "111111101110011010000111110" OR uut_a_1_0 /= "000000000000011101101110111" OR uut_a_1_1 /= "000000100111101110001111111" OR uut_a_1_2 /= "000000000101100100110011101" OR uut_a_1_3 /= "111111111111110000010101010" OR uut_a_1_4 /= "111111101011000100011010000" OR uut_a_1_5 /= "111111111101000011111111001" OR uut_a_2_0 /= "000000000000000100001011000" OR uut_a_2_1 /= "000000000101100100110011101" OR uut_a_2_2 /= "000000000000110010000101000" OR uut_a_2_3 /= "111111111111111101110011010" OR uut_a_2_4 /= "111111111101000011111111001" OR uut_a_2_5 /= "111111111111100101100111001" OR uut_a_3_0 /= "111111111110100010001011010" OR uut_a_3_1 /= "111110000010101010000111001" OR uut_a_3_2 /= "111111101110011010000111110" OR uut_a_3_3 /= "000000000000110001011100000" OR uut_a_3_4 /= "000001000010000010111111010" OR uut_a_3_5 /= "000000001001010001010000110" OR uut_a_4_0 /= "111111111111110000010101010" OR uut_a_4_1 /= "111111101011000100011010000" OR uut_a_4_2 /= "111111111101000011111111001" OR uut_a_4_3 /= "000000000000001000010000010" OR uut_a_4_4 /= "000000001011000001110111111" OR uut_a_4_5 /= "000000000001100011000100011" OR uut_a_5_0 /= "111111111111111101110011010" OR uut_a_5_1 /= "111111111101000011111111001" OR uut_a_5_2 /= "111111111111100101100111001" OR uut_a_5_3 /= "000000000000000001001010001" OR uut_a_5_4 /= "000000000001100011000100011" OR uut_a_5_5 /= "000000000000001101111001111" THEN
              FAIL <= '1';
              FAIL_NUM <= "01100001";
              state <= "11111101";
            ELSE
              state <= "01101111";
            END IF;
            uut_rst <= '0';
          WHEN "01101111" =>
            uut_coord_shift <= "1010";
            uut_x <= "001110110000";
            uut_y <= "001001010111";
            uut_fx <= "0101010101";
            uut_fy <= "1110011000";
            uut_ft <= "0100000000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000011000000100100" OR uut_a_0_1 /= "111111001000001001011010011" OR uut_a_0_2 /= "000010110101011110011001011" OR uut_a_0_3 /= "111111111111000011010010010" OR uut_a_0_4 /= "000010001100111000001001111" OR uut_a_0_5 /= "111000110110010001000101101" OR uut_a_1_0 /= "111111111111111001000001001" OR uut_a_1_1 /= "000000010000001100110001010" OR uut_a_1_2 /= "111111001011010111010111110" OR uut_a_1_3 /= "000000000000010001100111000" OR uut_a_1_4 /= "111111010111001000111101101" OR uut_a_1_5 /= "000010000100110000101010110" OR uut_a_2_0 /= "000000000000010110101011110" OR uut_a_2_1 /= "111111001011010111010111110" OR uut_a_2_2 /= "000010101011000001001101010" OR uut_a_2_3 /= "111111111111000110110010001" OR uut_a_2_4 /= "000010000100110000101010110" OR uut_a_2_5 /= "111001010000101000111110100" OR uut_a_3_0 /= "111111111111000011010010010" OR uut_a_3_1 /= "000010001100111000001001111" OR uut_a_3_2 /= "111000110110010001000101101" OR uut_a_3_3 /= "000000000010011001001001000" OR uut_a_3_4 /= "111010011100101010100111100" OR uut_a_3_5 /= "010010000010100010010110100" OR uut_a_4_0 /= "000000000000010001100111000" OR uut_a_4_1 /= "111111010111001000111101101" OR uut_a_4_2 /= "000010000100110000101010110" OR uut_a_4_3 /= "111111111111010011100101010" OR uut_a_4_4 /= "000001100111000011111000111" OR uut_a_4_5 /= "111010110001001000111010010" OR uut_a_5_0 /= "111111111111000110110010001" OR uut_a_5_1 /= "000010000100110000101010110" OR uut_a_5_2 /= "111001010000101000111110100" OR uut_a_5_3 /= "000000000010010000010100010" OR uut_a_5_4 /= "111010110001001000111010010" OR uut_a_5_5 /= "010001000000000000111111110" THEN
              FAIL <= '1';
              FAIL_NUM <= "01100010";
              state <= "11111101";
            ELSE
              state <= "01110000";
            END IF;
            uut_rst <= '0';
          WHEN "01110000" =>
            uut_coord_shift <= "1010";
            uut_x <= "010101011101";
            uut_y <= "110100101001";
            uut_fx <= "0000110110";
            uut_fy <= "0111101011";
            uut_ft <= "0000110010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000010001111010000000" OR uut_a_0_1 /= "111100111001111010010010011" OR uut_a_0_2 /= "110101111001001000011101111" OR uut_a_0_3 /= "000000000001001001010011110" OR uut_a_0_4 /= "111110011010101000001100001" OR uut_a_0_5 /= "111010110100111101110100010" OR uut_a_1_0 /= "111111111111100111001111010" OR uut_a_1_1 /= "000000100010001111010111001" OR uut_a_1_2 /= "000001101111110011111110010" OR uut_a_1_3 /= "111111111111110011010101000" OR uut_a_1_4 /= "000000010001100001011011011" OR uut_a_1_5 /= "000000111001001110000100001" OR uut_a_2_0 /= "111111111110101111001001000" OR uut_a_2_1 /= "000001101111110011111110010" OR uut_a_2_2 /= "000101101101001000000110000" OR uut_a_2_3 /= "111111111111010110100111101" OR uut_a_2_4 /= "000000111001001110000100001" OR uut_a_2_5 /= "000010111010110110100110111" OR uut_a_3_0 /= "000000000001001001010011110" OR uut_a_3_1 /= "111110011010101000001100001" OR uut_a_3_2 /= "111010110100111101110100010" OR uut_a_3_3 /= "000000000000100101100001000" OR uut_a_3_4 /= "111111001100000111110111100" OR uut_a_3_5 /= "111101010110100101111111000" OR uut_a_4_0 /= "111111111111110011010101000" OR uut_a_4_1 /= "000000010001100001011011011" OR uut_a_4_2 /= "000000111001001110000100001" OR uut_a_4_3 /= "111111111111111001100000111" OR uut_a_4_4 /= "000000001000111101111000111" OR uut_a_4_5 /= "000000011101010010000011110" OR uut_a_5_0 /= "111111111111010110100111101" OR uut_a_5_1 /= "000000111001001110000100001" OR uut_a_5_2 /= "000010111010110110100110111" OR uut_a_5_3 /= "111111111111101010110100101" OR uut_a_5_4 /= "000000011101010010000011110" OR uut_a_5_5 /= "000001011111100111110011110" THEN
              FAIL <= '1';
              FAIL_NUM <= "01100011";
              state <= "11111101";
            ELSE
              state <= "01110001";
            END IF;
            uut_rst <= '0';
          WHEN "01110001" =>
            uut_coord_shift <= "1010";
            uut_x <= "110101001010";
            uut_y <= "000111101001";
            uut_fx <= "1101110001";
            uut_fy <= "0100000111";
            uut_ft <= "1110101000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001111011000011001" OR uut_a_0_1 /= "010001011001001101010001011" OR uut_a_0_2 /= "001011111010010100110111000" OR uut_a_0_3 /= "111111111110101001111101101" OR uut_a_0_4 /= "110011110101101001000101000" OR uut_a_0_5 /= "110111101010111110101011000" OR uut_a_1_0 /= "000000000001000101100100110" OR uut_a_1_1 /= "001001110101011100001100010" OR uut_a_1_2 /= "000110101111000010101010111" OR uut_a_1_3 /= "111111111111001111010110100" OR uut_a_1_4 /= "111001000111111001001010100" OR uut_a_1_5 /= "111011010010100111010011111" OR uut_a_2_0 /= "000000000000101111101001010" OR uut_a_2_1 /= "000110101111000010101010111" OR uut_a_2_2 /= "000100100111001011011000111" OR uut_a_2_3 /= "111111111111011110101011111" OR uut_a_2_4 /= "111011010010100111010011111" OR uut_a_2_5 /= "111100110001100111000101000" OR uut_a_3_0 /= "111111111110101001111101101" OR uut_a_3_1 /= "110011110101101001000101000" OR uut_a_3_2 /= "110111101010111110101011000" OR uut_a_3_3 /= "000000000000111100001010000" OR uut_a_3_4 /= "001000100000001110110000000" OR uut_a_3_5 /= "000101110100101100001001011" OR uut_a_4_0 /= "111111111111001111010110100" OR uut_a_4_1 /= "111001000111111001001010100" OR uut_a_4_2 /= "111011010010100111010011111" OR uut_a_4_3 /= "000000000000100010000000111" OR uut_a_4_4 /= "000100110011101110010101110" OR uut_a_4_5 /= "000011010010101110101101100" OR uut_a_5_0 /= "111111111111011110101011111" OR uut_a_5_1 /= "111011010010100111010011111" OR uut_a_5_2 /= "111100110001100111000101000" OR uut_a_5_3 /= "000000000000010111010010110" OR uut_a_5_4 /= "000011010010101110101101100" OR uut_a_5_5 /= "000010010000010011101110000" THEN
              FAIL <= '1';
              FAIL_NUM <= "01100100";
              state <= "11111101";
            ELSE
              state <= "01110010";
            END IF;
            uut_rst <= '0';
          WHEN "01110010" =>
            uut_coord_shift <= "1010";
            uut_x <= "111111100001";
            uut_y <= "001100011101";
            uut_fx <= "0111100100";
            uut_fy <= "1101010000";
            uut_ft <= "0101011010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000111101000010" OR uut_a_0_1 /= "000001000010000110011111111" OR uut_a_0_2 /= "111110010000010111000100100" OR uut_a_0_3 /= "111111111111110011001111100" OR uut_a_0_4 /= "111110010001011110100110101" OR uut_a_0_5 /= "000010111010101010010100011" OR uut_a_1_0 /= "000000000000000100001000011" OR uut_a_1_1 /= "000000100011110010110101001" OR uut_a_1_2 /= "111111000011100010111111100" OR uut_a_1_3 /= "111111111111111001000101111" OR uut_a_1_4 /= "111111000100001001101110101" OR uut_a_1_5 /= "000001100101000100111110101" OR uut_a_2_0 /= "111111111111111001000001011" OR uut_a_2_1 /= "111111000011100010111111100" OR uut_a_2_2 /= "000001100110000110011001100" OR uut_a_2_3 /= "000000000000001011101010101" OR uut_a_2_4 /= "000001100101000100111110101" OR uut_a_2_5 /= "111101010101010010011110111" OR uut_a_3_0 /= "111111111111110011001111100" OR uut_a_3_1 /= "111110010001011110100110101" OR uut_a_3_2 /= "000010111010101010010100011" OR uut_a_3_3 /= "000000000000010101010101000" OR uut_a_3_4 /= "000010111000110010101101110" OR uut_a_3_5 /= "111011000111111001110000001" OR uut_a_4_0 /= "111111111111111001000101111" OR uut_a_4_1 /= "111111000100001001101110101" OR uut_a_4_2 /= "000001100101000100111110101" OR uut_a_4_3 /= "000000000000001011100011001" OR uut_a_4_4 /= "000001100100000100001101101" OR uut_a_4_5 /= "111101010110111111110111100" OR uut_a_5_0 /= "000000000000001011101010101" OR uut_a_5_1 /= "000001100101000100111110101" OR uut_a_5_2 /= "111101010101010010011110111" OR uut_a_5_3 /= "111111111111101100011111100" OR uut_a_5_4 /= "111101010110111111110111100" OR uut_a_5_5 /= "000100011101011011011101100" THEN
              FAIL <= '1';
              FAIL_NUM <= "01100101";
              state <= "11111101";
            ELSE
              state <= "01110011";
            END IF;
            uut_rst <= '0';
          WHEN "01110011" =>
            uut_coord_shift <= "1010";
            uut_x <= "001111010011";
            uut_y <= "011101000100";
            uut_fx <= "1000100001";
            uut_fy <= "1101101101";
            uut_ft <= "0010100111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000001111010011000" OR uut_a_0_1 /= "111101111001000100101000110" OR uut_a_0_2 /= "111110001111000011111111101" OR uut_a_0_3 /= "111111111111111110000000110" OR uut_a_0_4 /= "000000010001100010000110111" OR uut_a_0_5 /= "000000001110101011001110110" OR uut_a_1_0 /= "111111111111110111100100010" OR uut_a_1_1 /= "000001001010011000011010010" OR uut_a_1_2 /= "000000111110010000100101000" OR uut_a_1_3 /= "000000000000000001000110001" OR uut_a_1_4 /= "111111110110010101011010100" OR uut_a_1_5 /= "111111110111111010001110101" OR uut_a_2_0 /= "111111111111111000111100001" OR uut_a_2_1 /= "000000111110010000100101000" OR uut_a_2_2 /= "000000110100000111001011111" OR uut_a_2_3 /= "000000000000000000111010101" OR uut_a_2_4 /= "111111110111111010001110101" OR uut_a_2_5 /= "111111111001001110100111010" OR uut_a_3_0 /= "111111111111111110000000110" OR uut_a_3_1 /= "000000010001100010000110111" OR uut_a_3_2 /= "000000001110101011001110110" OR uut_a_3_3 /= "000000000000000000010000100" OR uut_a_3_4 /= "111111111101101110001100000" OR uut_a_3_5 /= "111111111110000101111100111" OR uut_a_4_0 /= "000000000000000001000110001" OR uut_a_4_1 /= "111111110110010101011010100" OR uut_a_4_2 /= "111111110111111010001110101" OR uut_a_4_3 /= "111111111111111111110110111" OR uut_a_4_4 /= "000000000001010000011000011" OR uut_a_4_5 /= "000000000001000011010001111" OR uut_a_5_0 /= "000000000000000000111010101" OR uut_a_5_1 /= "111111110111111010001110101" OR uut_a_5_2 /= "111111111001001110100111010" OR uut_a_5_3 /= "111111111111111111111000010" OR uut_a_5_4 /= "000000000001000011010001111" OR uut_a_5_5 /= "000000000000111000010100001" THEN
              FAIL <= '1';
              FAIL_NUM <= "01100110";
              state <= "11111101";
            ELSE
              state <= "01110100";
            END IF;
            uut_rst <= '0';
          WHEN "01110100" =>
            uut_coord_shift <= "1010";
            uut_x <= "110010000010";
            uut_y <= "101110110000";
            uut_fx <= "0011011000";
            uut_fy <= "0010000000";
            uut_ft <= "0001011101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000110111110010001" OR uut_a_0_1 /= "111000101001110000111101100" OR uut_a_0_2 /= "110110111111110111010011011" OR uut_a_0_3 /= "000000000000101101000011100" OR uut_a_0_4 /= "111010000100001100011110000" OR uut_a_0_5 /= "111000101110101010001101001" OR uut_a_1_0 /= "111111111111100010100111000" OR uut_a_1_1 /= "000011110111101111101111000" OR uut_a_1_2 /= "000100101111100010100101010" OR uut_a_1_3 /= "111111111111101000010000110" OR uut_a_1_4 /= "000011001000000110100011100" OR uut_a_1_5 /= "000011110101001010101100110" OR uut_a_2_0 /= "111111111111011011111111011" OR uut_a_2_1 /= "000100101111100010100101010" OR uut_a_2_2 /= "000101110011111001100111010" OR uut_a_2_3 /= "111111111111100010111010101" OR uut_a_2_4 /= "000011110101001010101100110" OR uut_a_2_5 /= "000100101100011000011000010" OR uut_a_3_0 /= "000000000000101101000011100" OR uut_a_3_1 /= "111010000100001100011110000" OR uut_a_3_2 /= "111000101110101010001101001" OR uut_a_3_3 /= "000000000000100100011001000" OR uut_a_3_4 /= "111011001101001110111111101" OR uut_a_3_5 /= "111010001000001001011110010" OR uut_a_4_0 /= "111111111111101000010000110" OR uut_a_4_1 /= "000011001000000110100011100" OR uut_a_4_2 /= "000011110101001010101100110" OR uut_a_4_3 /= "111111111111101100110100111" OR uut_a_4_4 /= "000010100001100111110000011" OR uut_a_4_5 /= "000011000110000001010000100" OR uut_a_5_0 /= "111111111111100010111010101" OR uut_a_5_1 /= "000011110101001010101100110" OR uut_a_5_2 /= "000100101100011000011000010" OR uut_a_5_3 /= "111111111111101000100000100" OR uut_a_5_4 /= "000011000110000001010000100" OR uut_a_5_5 /= "000011110010100111011000100" THEN
              FAIL <= '1';
              FAIL_NUM <= "01100111";
              state <= "11111101";
            ELSE
              state <= "01110101";
            END IF;
            uut_rst <= '0';
          WHEN "01110101" =>
            uut_coord_shift <= "1010";
            uut_x <= "001010010001";
            uut_y <= "100011000011";
            uut_fx <= "1101100101";
            uut_fy <= "1111001110";
            uut_ft <= "1011110111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001010010011110110" OR uut_a_0_1 /= "101111110101000111110010101" OR uut_a_0_2 /= "110010111001101010001000110" OR uut_a_0_3 /= "000000000000000010000000011" OR uut_a_0_4 /= "111111100110110100100000101" OR uut_a_0_5 /= "111111101011100110100011011" OR uut_a_1_0 /= "111111111110111111010100011" OR uut_a_1_1 /= "001100101011100001111100111" OR uut_a_1_2 /= "001010010001011010010001001" OR uut_a_1_3 /= "111111111111111110011011010" OR uut_a_1_4 /= "000000010011101111101100100" OR uut_a_1_5 /= "000000001111111111101101000" OR uut_a_2_0 /= "111111111111001011100110101" OR uut_a_2_1 /= "001010010001011010010001001" OR uut_a_2_2 /= "001000010100100011110100110" OR uut_a_2_3 /= "111111111111111110101110011" OR uut_a_2_4 /= "000000001111111111101101000" OR uut_a_2_5 /= "000000001100111101010010100" OR uut_a_3_0 /= "000000000000000010000000011" OR uut_a_3_1 /= "111111100110110100100000101" OR uut_a_3_2 /= "111111101011100110100011011" OR uut_a_3_3 /= "000000000000000000000011001" OR uut_a_3_4 /= "111111111111011000110010101" OR uut_a_3_5 /= "111111111111100000001111001" OR uut_a_4_0 /= "111111111111111110011011010" OR uut_a_4_1 /= "000000010011101111101100100" OR uut_a_4_2 /= "000000001111111111101101000" OR uut_a_4_3 /= "111111111111111111111101100" OR uut_a_4_4 /= "000000000000011110101111110" OR uut_a_4_5 /= "000000000000011000111010000" OR uut_a_5_0 /= "111111111111111110101110011" OR uut_a_5_1 /= "000000001111111111101101000" OR uut_a_5_2 /= "000000001100111101010010100" OR uut_a_5_3 /= "111111111111111111111110000" OR uut_a_5_4 /= "000000000000011000111010000" OR uut_a_5_5 /= "000000000000010100001011010" THEN
              FAIL <= '1';
              FAIL_NUM <= "01101000";
              state <= "11111101";
            ELSE
              state <= "01110110";
            END IF;
            uut_rst <= '0';
          WHEN "01110110" =>
            uut_coord_shift <= "1010";
            uut_x <= "001101110000";
            uut_y <= "010110110010";
            uut_fx <= "1100100000";
            uut_fy <= "0011101101";
            uut_ft <= "1010001101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001101010011111010" OR uut_a_0_1 /= "010101000100100101001001011" OR uut_a_0_2 /= "101010101001111100101110000" OR uut_a_0_3 /= "111111111111110010100010111" OR uut_a_0_4 /= "111101010101100111110110001" OR uut_a_0_5 /= "000010101100100101011010101" OR uut_a_1_0 /= "000000000001010100010010010" OR uut_a_1_1 /= "010000101011011010000001110" OR uut_a_1_2 /= "101111000110110000111101110" OR uut_a_1_3 /= "111111111111110101010110011" OR uut_a_1_4 /= "111101111001001001010100011" OR uut_a_1_5 /= "000010001000100110011111011" OR uut_a_2_0 /= "111111111110101010100111110" OR uut_a_2_1 /= "101111000110110000111101110" OR uut_a_2_2 /= "010001000111001111100000010" OR uut_a_2_3 /= "000000000000001010110010010" OR uut_a_2_4 /= "000010001000100110011111011" OR uut_a_2_5 /= "111101110101101000010000000" OR uut_a_3_0 /= "111111111111110010100010111" OR uut_a_3_1 /= "111101010101100111110110001" OR uut_a_3_2 /= "000010101100100101011010101" OR uut_a_3_3 /= "000000000000000001101100110" OR uut_a_3_4 /= "000000010101100001100111001" OR uut_a_3_5 /= "111111101010001100100010100" OR uut_a_4_0 /= "111111111111110101010110011" OR uut_a_4_1 /= "111101111001001001010100011" OR uut_a_4_2 /= "000010001000100110011111011" OR uut_a_4_3 /= "000000000000000001010110000" OR uut_a_4_4 /= "000000010001000010011000101" OR uut_a_4_5 /= "111111101110101111011111010" OR uut_a_5_0 /= "000000000000001010110010010" OR uut_a_5_1 /= "000010001000100110011111011" OR uut_a_5_2 /= "111101110101101000010000000" OR uut_a_5_3 /= "111111111111111110101000110" OR uut_a_5_4 /= "111111101110101111011111010" OR uut_a_5_5 /= "000000010001011110110100100" THEN
              FAIL <= '1';
              FAIL_NUM <= "01101001";
              state <= "11111101";
            ELSE
              state <= "01110111";
            END IF;
            uut_rst <= '0';
          WHEN "01110111" =>
            uut_coord_shift <= "1010";
            uut_x <= "010101100011";
            uut_y <= "101000111000";
            uut_fx <= "0001011010";
            uut_fy <= "1101110111";
            uut_ft <= "0100111010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000001101010010110" OR uut_a_0_1 /= "111110110000000010000001001" OR uut_a_0_2 /= "111101110111100010001100101" OR uut_a_0_3 /= "000000000000010111111011011" OR uut_a_0_4 /= "111101110000000011101000100" OR uut_a_0_5 /= "111100001010010111001010000" OR uut_a_1_0 /= "111111111111111011000000001" OR uut_a_1_1 /= "000000011110000100001111011" OR uut_a_1_2 /= "000000110011010011101101000" OR uut_a_1_3 /= "111111111111110111000000001" OR uut_a_1_4 /= "000000110110000111101000100" OR uut_a_1_5 /= "000001011100010110101010110" OR uut_a_2_0 /= "111111111111110111011110001" OR uut_a_2_1 /= "000000110011010011101101000" OR uut_a_2_2 /= "000001010111100011100111101" OR uut_a_2_3 /= "111111111111110000101001011" OR uut_a_2_4 /= "000001011100010110101010110" OR uut_a_2_5 /= "000010011101100110100001000" OR uut_a_3_0 /= "000000000000010111111011011" OR uut_a_3_1 /= "111101110000000011101000100" OR uut_a_3_2 /= "111100001010010111001010000" OR uut_a_3_3 /= "000000000000101011000100100" OR uut_a_3_4 /= "111011111100111001101111011" OR uut_a_3_5 /= "111001000101110110011110111" OR uut_a_4_0 /= "111111111111110111000000001" OR uut_a_4_1 /= "000000110110000111101000100" OR uut_a_4_2 /= "000001011100010110101010110" OR uut_a_4_3 /= "111111111111101111110011100" OR uut_a_4_4 /= "000001100001011010100010100" OR uut_a_4_5 /= "000010100110001111001100111" OR uut_a_5_0 /= "111111111111110000101001011" OR uut_a_5_1 /= "000001011100010110101010110" OR uut_a_5_2 /= "000010011101100110100001000" OR uut_a_5_3 /= "111111111111100100010111011" OR uut_a_5_4 /= "000010100110001111001100111" OR uut_a_5_5 /= "000100011011101011101110110" THEN
              FAIL <= '1';
              FAIL_NUM <= "01101010";
              state <= "11111101";
            ELSE
              state <= "01111000";
            END IF;
            uut_rst <= '0';
          WHEN "01111000" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000000000";
            uut_y <= "111111111111";
            uut_fx <= "0110000010";
            uut_fy <= "1101101010";
            uut_ft <= "1111001100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001010001010010000" OR uut_a_0_1 /= "010000100000101010000000000" OR uut_a_0_2 /= "000101001111010010010000000" OR uut_a_0_3 /= "000000000000010110010100000" OR uut_a_0_4 /= "000100100010000100000000000" OR uut_a_0_5 /= "000001011100000010100000000" OR uut_a_1_0 /= "000000000001000010000010101" OR uut_a_1_1 /= "001101011010100010001000000" OR uut_a_1_2 /= "000100010000011010110101000" OR uut_a_1_3 /= "000000000000010010001000010" OR uut_a_1_4 /= "000011101011101011010000000" OR uut_a_1_5 /= "000001001010110010000010000" OR uut_a_2_0 /= "000000000000010100111101001" OR uut_a_2_1 /= "000100010000011010110101000" OR uut_a_2_2 /= "000001010110011100001101001" OR uut_a_2_3 /= "000000000000000101110000001" OR uut_a_2_4 /= "000001001010110010000010000" OR uut_a_2_5 /= "000000010111101110101001010" OR uut_a_3_0 /= "000000000000010110010100000" OR uut_a_3_1 /= "000100100010000100000000000" OR uut_a_3_2 /= "000001011100000010100000000" OR uut_a_3_3 /= "000000000000000110001000000" OR uut_a_3_4 /= "000001001111101000000000000" OR uut_a_3_5 /= "000000011001010001000000000" OR uut_a_4_0 /= "000000000000010010001000010" OR uut_a_4_1 /= "000011101011101011010000000" OR uut_a_4_2 /= "000001001010110010000010000" OR uut_a_4_3 /= "000000000000000100111110100" OR uut_a_4_4 /= "000001000000101100100000000" OR uut_a_4_5 /= "000000010100100001110100000" OR uut_a_5_0 /= "000000000000000101110000001" OR uut_a_5_1 /= "000001001010110010000010000" OR uut_a_5_2 /= "000000010111101110101001010" OR uut_a_5_3 /= "000000000000000001100101000" OR uut_a_5_4 /= "000000010100100001110100000" OR uut_a_5_5 /= "000000000110100000111000100" THEN
              FAIL <= '1';
              FAIL_NUM <= "01101011";
              state <= "11111101";
            ELSE
              state <= "01111001";
            END IF;
            uut_rst <= '0';
          WHEN "01111001" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000111011";
            uut_y <= "111111000110";
            uut_fx <= "0111100100";
            uut_fy <= "1011000010";
            uut_ft <= "0010101011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001111111000000001" OR uut_a_0_1 /= "000000000100111101100000010" OR uut_a_0_2 /= "111011101011001011001110100" OR uut_a_0_3 /= "000000000001001111011100000" OR uut_a_0_4 /= "000000000011000110100110001" OR uut_a_0_5 /= "111101010010110110010101010" OR uut_a_1_0 /= "000000000000000000010011110" OR uut_a_1_1 /= "000000000000000000110001100" OR uut_a_1_2 /= "111111111111010100101111110" OR uut_a_1_3 /= "000000000000000000001100011" OR uut_a_1_4 /= "000000000000000000011111000" OR uut_a_1_5 /= "111111111111100100111100011" OR uut_a_2_0 /= "111111111111101110101100101" OR uut_a_2_1 /= "111111111111010100101111110" OR uut_a_2_2 /= "000000100101101101100100000" OR uut_a_2_3 /= "111111111111110101001011011" OR uut_a_2_4 /= "111111111111100100111100011" OR uut_a_2_5 /= "000000010111100101101010010" OR uut_a_3_0 /= "000000000001001111011100000" OR uut_a_3_1 /= "000000000011000110100110001" OR uut_a_3_2 /= "111101010010110110010101010" OR uut_a_3_3 /= "000000000000110001101100000" OR uut_a_3_4 /= "000000000001111100001110000" OR uut_a_3_5 /= "111110010011101100100001101" OR uut_a_4_0 /= "000000000000000000001100011" OR uut_a_4_1 /= "000000000000000000011111000" OR uut_a_4_2 /= "111111111111100100111100011" OR uut_a_4_3 /= "000000000000000000000111110" OR uut_a_4_4 /= "000000000000000000010011011" OR uut_a_4_5 /= "111111111111101111000100111" OR uut_a_5_0 /= "111111111111110101001011011" OR uut_a_5_1 /= "111111111111100100111100011" OR uut_a_5_2 /= "000000010111100101101010010" OR uut_a_5_3 /= "111111111111111001001110110" OR uut_a_5_4 /= "111111111111101111000100111" OR uut_a_5_5 /= "000000001110110000010001110" THEN
              FAIL <= '1';
              FAIL_NUM <= "01101100";
              state <= "11111101";
            ELSE
              state <= "01111010";
            END IF;
            uut_rst <= '0';
          WHEN "01111010" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000001011";
            uut_y <= "000000010110";
            uut_fx <= "1101110010";
            uut_fy <= "0001111011";
            uut_ft <= "0100111111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000110001111000" OR uut_a_0_1 /= "000001001110101010101001101" OR uut_a_0_2 /= "111110110111101101101110110" OR uut_a_0_3 /= "111111111111100111110101010" OR uut_a_0_4 /= "111011001111000101001001110" OR uut_a_0_5 /= "000100011000001011111010001" OR uut_a_1_0 /= "000000000000000100111010101" OR uut_a_1_1 /= "000000111110000010001100100" OR uut_a_1_2 /= "111111000110111111110110000" OR uut_a_1_3 /= "111111111111101100111100010" OR uut_a_1_4 /= "111100001111100011000110000" OR uut_a_1_5 /= "000011011100111100101000111" OR uut_a_2_0 /= "111111111111111011011110110" OR uut_a_2_1 /= "111111000110111111110110000" OR uut_a_2_2 /= "000000110100011000001111001" OR uut_a_2_3 /= "000000000000010001100000101" OR uut_a_2_4 /= "000011011100111100101000111" OR uut_a_2_5 /= "111100110100111110010111110" OR uut_a_3_0 /= "111111111111100111110101010" OR uut_a_3_1 /= "111011001111000101001001110" OR uut_a_3_2 /= "000100011000001011111010001" OR uut_a_3_3 /= "000000000001011101101011001" OR uut_a_3_4 /= "010010011101111001100111011" OR uut_a_3_5 /= "101111000001111110000001010" OR uut_a_4_0 /= "111111111111101100111100010" OR uut_a_4_1 /= "111100001111100011000110000" OR uut_a_4_2 /= "000011011100111100101000111" OR uut_a_4_3 /= "000000000001001001110111100" OR uut_a_4_4 /= "001110100100000001000001110" OR uut_a_4_5 /= "110010100111100101011000000" OR uut_a_5_0 /= "000000000000010001100000101" OR uut_a_5_1 /= "000011011100111100101000111" OR uut_a_5_2 /= "111100110100111110010111110" OR uut_a_5_3 /= "111111111110111100000111111" OR uut_a_5_4 /= "110010100111100101011000000" OR uut_a_5_5 /= "001100010010111100101011110" THEN
              FAIL <= '1';
              FAIL_NUM <= "01101101";
              state <= "11111101";
            ELSE
              state <= "01111011";
            END IF;
            uut_rst <= '0';
          WHEN "01111011" =>
            uut_coord_shift <= "0101";
            uut_x <= "111111000011";
            uut_y <= "111111001011";
            uut_fx <= "0111100110";
            uut_fy <= "0010011011";
            uut_ft <= "1011101101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000001100100000000" OR uut_a_0_1 /= "000001010101010110100000000" OR uut_a_0_2 /= "000000101111010001000000000" OR uut_a_0_3 /= "111111111111011101001010000" OR uut_a_0_4 /= "111100010010000101010010000" OR uut_a_0_5 /= "111101111100001111110100000" OR uut_a_1_0 /= "000000000000000101010101011" OR uut_a_1_1 /= "000000100100011011001010100" OR uut_a_1_2 /= "000000010100001010111100010" OR uut_a_1_3 /= "111111111111110001001000010" OR uut_a_1_4 /= "111110011010011101111000001" OR uut_a_1_5 /= "111111000111110001011111111" OR uut_a_2_0 /= "000000000000000010111101000" OR uut_a_2_1 /= "000000010100001010111100010" OR uut_a_2_2 /= "000000001011001010111001001" OR uut_a_2_3 /= "111111111111110111110000111" OR uut_a_2_4 /= "111111000111110001011111111" OR uut_a_2_5 /= "111111100000110111001111001" OR uut_a_3_0 /= "111111111111011101001010000" OR uut_a_3_1 /= "111100010010000101010010000" OR uut_a_3_2 /= "111101111100001111110100000" OR uut_a_3_3 /= "000000000001100001001000001" OR uut_a_3_4 /= "001010010111001100011110101" OR uut_a_3_5 /= "000101101111010000101110010" OR uut_a_4_0 /= "111111111111110001001000010" OR uut_a_4_1 /= "111110011010011101111000001" OR uut_a_4_2 /= "111111000111110001011111111" OR uut_a_4_3 /= "000000000000101001011100110" OR uut_a_4_4 /= "000100011011000001100000110" OR uut_a_4_5 /= "000010011100101110110100101" OR uut_a_5_0 /= "111111111111110111110000111" OR uut_a_5_1 /= "111111000111110001011111111" OR uut_a_5_2 /= "111111100000110111001111001" OR uut_a_5_3 /= "000000000000010110111101000" OR uut_a_5_4 /= "000010011100101110110100101" OR uut_a_5_5 /= "000001010110110010110100111" THEN
              FAIL <= '1';
              FAIL_NUM <= "01101110";
              state <= "11111101";
            ELSE
              state <= "01111100";
            END IF;
            uut_rst <= '0';
          WHEN "01111100" =>
            uut_coord_shift <= "0101";
            uut_x <= "111111110100";
            uut_y <= "111111010000";
            uut_fx <= "1100010011";
            uut_fy <= "1100001000";
            uut_ft <= "1101010100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000111000110001110" OR uut_a_0_1 /= "000110100010101111001000110" OR uut_a_0_2 /= "000100001001101100111101011" OR uut_a_0_3 /= "111111111111101110101011110" OR uut_a_0_4 /= "111110000000010010101010000" OR uut_a_0_5 /= "111110101110111101101111001" OR uut_a_1_0 /= "000000000000011010001010111" OR uut_a_1_1 /= "000011000001000000101110100" OR uut_a_1_2 /= "000001111010011110001110010" OR uut_a_1_3 /= "111111111111111000000001001" OR uut_a_1_4 /= "111111000101001000100110010" OR uut_a_1_5 /= "111111011010101001011101001" OR uut_a_2_0 /= "000000000000010000100110110" OR uut_a_2_1 /= "000001111010011110001110010" OR uut_a_2_2 /= "000001001101101101100111100" OR uut_a_2_3 /= "111111111111111010111011110" OR uut_a_2_4 /= "111111011010101001011101001" OR uut_a_2_5 /= "111111101000010011000111101" OR uut_a_3_0 /= "111111111111101110101011110" OR uut_a_3_1 /= "111110000000010010101010000" OR uut_a_3_2 /= "111110101110111101101111001" OR uut_a_3_3 /= "000000000000000101010010000" OR uut_a_3_4 /= "000000100110111100110000000" OR uut_a_3_5 /= "000000011000101101101111000" OR uut_a_4_0 /= "111111111111111000000001001" OR uut_a_4_1 /= "111111000101001000100110010" OR uut_a_4_2 /= "111111011010101001011101001" OR uut_a_4_3 /= "000000000000000010011011110" OR uut_a_4_4 /= "000000010001111101000000001" OR uut_a_4_5 /= "000000001011011001000101001" OR uut_a_5_0 /= "111111111111111010111011110" OR uut_a_5_1 /= "111111011010101001011101001" OR uut_a_5_2 /= "111111101000010011000111101" OR uut_a_5_3 /= "000000000000000001100010110" OR uut_a_5_4 /= "000000001011011001000101001" OR uut_a_5_5 /= "000000000111001110101000000" THEN
              FAIL <= '1';
              FAIL_NUM <= "01101111";
              state <= "11111101";
            ELSE
              state <= "01111101";
            END IF;
            uut_rst <= '0';
          WHEN "01111101" =>
            uut_coord_shift <= "0101";
            uut_x <= "111111010100";
            uut_y <= "111111101101";
            uut_fx <= "1001111101";
            uut_fy <= "0110001001";
            uut_ft <= "1001100001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000001011011001" OR uut_a_0_1 /= "000000001111010001011101010" OR uut_a_0_2 /= "111111110111111010011100000" OR uut_a_0_3 /= "000000000000001100111100100" OR uut_a_0_4 /= "000010001010110111101000001" OR uut_a_0_5 /= "111110110110011110000001100" OR uut_a_1_0 /= "000000000000000000111101000" OR uut_a_1_1 /= "000000001010001111010011000" OR uut_a_1_2 /= "111111111010100101000001011" OR uut_a_1_3 /= "000000000000001000101011011" OR uut_a_1_4 /= "000001011101000110010110110" OR uut_a_1_5 /= "111111001110101101000100001" OR uut_a_2_0 /= "111111111111111111011111101" OR uut_a_2_1 /= "111111111010100101000001011" OR uut_a_2_2 /= "000000000010110111101110010" OR uut_a_2_3 /= "111111111111111011011001111" OR uut_a_2_4 /= "111111001110101101000100001" OR uut_a_2_5 /= "000000011010000110100001111" OR uut_a_3_0 /= "000000000000001100111100100" OR uut_a_3_1 /= "000010001010110111101000001" OR uut_a_3_2 /= "111110110110011110000001100" OR uut_a_3_3 /= "000000000001110101101101110" OR uut_a_3_4 /= "010011101110101011100100110" OR uut_a_3_5 /= "110101100011011010011110100" OR uut_a_4_0 /= "000000000000001000101011011" OR uut_a_4_1 /= "000001011101000110010110110" OR uut_a_4_2 /= "111111001110101101000100001" OR uut_a_4_3 /= "000000000001001110111010101" OR uut_a_4_4 /= "001101001110100000111001101" OR uut_a_4_5 /= "111000111111110001011110000" OR uut_a_5_0 /= "111111111111111011011001111" OR uut_a_5_1 /= "111111001110101101000100001" OR uut_a_5_2 /= "000000011010000110100001111" OR uut_a_5_3 /= "111111111111010110001101101" OR uut_a_5_4 /= "111000111111110001011110000" OR uut_a_5_5 /= "000011101101010101011100011" THEN
              FAIL <= '1';
              FAIL_NUM <= "01110000";
              state <= "11111101";
            ELSE
              state <= "01111110";
            END IF;
            uut_rst <= '0';
          WHEN "01111110" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000110111";
            uut_y <= "111111110100";
            uut_fx <= "1000110001";
            uut_fy <= "1101011111";
            uut_ft <= "0011110010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000001001111111000" OR uut_a_0_1 /= "111111001001110111010000001" OR uut_a_0_2 /= "000000100110001001010011001" OR uut_a_0_3 /= "111111111111101101101000101" OR uut_a_0_4 /= "000001100011100100001110100" OR uut_a_0_5 /= "111110111001110110000011101" OR uut_a_1_0 /= "111111111111111100100111011" OR uut_a_1_1 /= "000000010010010110000101101" OR uut_a_1_2 /= "111111110011000100101110010" OR uut_a_1_3 /= "000000000000000110001110010" OR uut_a_1_4 /= "111111011110010000101010010" OR uut_a_1_5 /= "000000010111110001011111100" OR uut_a_2_0 /= "000000000000000010011000100" OR uut_a_2_1 /= "111111110011000100101110010" OR uut_a_2_2 /= "000000001001000110111010000" OR uut_a_2_3 /= "111111111111111011100111011" OR uut_a_2_4 /= "000000010111110001011111100" OR uut_a_2_5 /= "111111101111001111111100000" OR uut_a_3_0 /= "111111111111101101101000101" OR uut_a_3_1 /= "000001100011100100001110100" OR uut_a_3_2 /= "111110111001110110000011101" OR uut_a_3_3 /= "000000000000100001110001100" OR uut_a_3_4 /= "111101001000111000011100101" OR uut_a_3_5 /= "000010000001000001101110011" OR uut_a_4_0 /= "000000000000000110001110010" OR uut_a_4_1 /= "111111011110010000101010010" OR uut_a_4_2 /= "000000010111110001011111100" OR uut_a_4_3 /= "111111111111110100100011100" OR uut_a_4_4 /= "000000111110000011010111110" OR uut_a_4_5 /= "111111010100010001101110100" OR uut_a_5_0 /= "111111111111111011100111011" OR uut_a_5_1 /= "000000010111110001011111100" OR uut_a_5_2 /= "111111101111001111111100000" OR uut_a_5_3 /= "000000000000001000000100000" OR uut_a_5_4 /= "111111010100010001101110100" OR uut_a_5_5 /= "000000011110110011101100010" THEN
              FAIL <= '1';
              FAIL_NUM <= "01110001";
              state <= "11111101";
            ELSE
              state <= "01111111";
            END IF;
            uut_rst <= '0';
          WHEN "01111111" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000100101";
            uut_y <= "000000000101";
            uut_fx <= "0010111111";
            uut_fy <= "0110010011";
            uut_ft <= "1000111000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001110010011000100" OR uut_a_0_1 /= "111111100100010011000100010" OR uut_a_0_2 /= "001011001000001101100011010" OR uut_a_0_3 /= "111111111111010110011010000" OR uut_a_0_4 /= "000000001010000100101101000" OR uut_a_0_5 /= "111011111101000000111001000" OR uut_a_1_0 /= "111111111111111110010001001" OR uut_a_1_1 /= "000000000000011010110101100" OR uut_a_1_2 /= "111111110101001110000010110" OR uut_a_1_3 /= "000000000000000000101000010" OR uut_a_1_4 /= "111111111111110110001111011" OR uut_a_1_5 /= "000000000011111010111001001" OR uut_a_2_0 /= "000000000000101100100000110" OR uut_a_2_1 /= "111111110101001110000010110" OR uut_a_2_2 /= "000100010101001010100001011" OR uut_a_2_3 /= "111111111111101111110100000" OR uut_a_2_4 /= "000000000011111010111001001" OR uut_a_2_5 /= "111110011011001101101000001" OR uut_a_3_0 /= "111111111111010110011010000" OR uut_a_3_1 /= "000000001010000100101101000" OR uut_a_3_2 /= "111011111101000000111001000" OR uut_a_3_3 /= "000000000000001111001000000" OR uut_a_3_4 /= "111111111100010101100100000" OR uut_a_3_5 /= "000001011110001011010100000" OR uut_a_4_0 /= "000000000000000000101000010" OR uut_a_4_1 /= "111111111111110110001111011" OR uut_a_4_2 /= "000000000011111010111001001" OR uut_a_4_3 /= "111111111111111111110001010" OR uut_a_4_4 /= "000000000000000011100011000" OR uut_a_4_5 /= "111111111110100100110001000" OR uut_a_5_0 /= "111111111111101111110100000" OR uut_a_5_1 /= "000000000011111010111001001" OR uut_a_5_2 /= "111110011011001101101000001" OR uut_a_5_3 /= "000000000000000101111000101" OR uut_a_5_4 /= "111111111110100100110001000" OR uut_a_5_5 /= "000000100100101001100101110" THEN
              FAIL <= '1';
              FAIL_NUM <= "01110010";
              state <= "11111101";
            ELSE
              state <= "10000000";
            END IF;
            uut_rst <= '0';
          WHEN "10000000" =>
            uut_coord_shift <= "0101";
            uut_x <= "111111100111";
            uut_y <= "111111000110";
            uut_fx <= "1011001000";
            uut_fy <= "0011100001";
            uut_ft <= "0011100011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001110000000010000" OR uut_a_0_1 /= "001101011000110111100010010" OR uut_a_0_2 /= "011001011011111101100001000" OR uut_a_0_3 /= "000000000000100010011000011" OR uut_a_0_4 /= "000100000110111101101010110" OR uut_a_0_5 /= "000111110011100110101001110" OR uut_a_1_0 /= "000000000000110101100011011" OR uut_a_1_1 /= "000110011001100110110011000" OR uut_a_1_2 /= "001100001010001101011100000" OR uut_a_1_3 /= "000000000000010000011011110" OR uut_a_1_4 /= "000001111101101101000010101" OR uut_a_1_5 /= "000011101110110100110000100" OR uut_a_2_0 /= "000000000001100101101111110" OR uut_a_2_1 /= "001100001010001101011100000" OR uut_a_2_2 /= "010111000110100001001111101" OR uut_a_2_3 /= "000000000000011111001110011" OR uut_a_2_4 /= "000011101110110100110000100" OR uut_a_2_5 /= "000111000101101111011110101" OR uut_a_3_0 /= "000000000000100010011000011" OR uut_a_3_1 /= "000100000110111101101010110" OR uut_a_3_2 /= "000111110011100110101001110" OR uut_a_3_3 /= "000000000000001010100011010" OR uut_a_3_4 /= "000001010000101100110110001" OR uut_a_3_5 /= "000010011001010100101011100" OR uut_a_4_0 /= "000000000000010000011011110" OR uut_a_4_1 /= "000001111101101101000010101" OR uut_a_4_2 /= "000011101110110100110000100" OR uut_a_4_3 /= "000000000000000101000010110" OR uut_a_4_4 /= "000000100110100100111100000" OR uut_a_4_5 /= "000001001001010010101110101" OR uut_a_5_0 /= "000000000000011111001110011" OR uut_a_5_1 /= "000011101110110100110000100" OR uut_a_5_2 /= "000111000101101111011110101" OR uut_a_5_3 /= "000000000000001001100101010" OR uut_a_5_4 /= "000001001001010010101110101" OR uut_a_5_5 /= "000010001011001111111010000" THEN
              FAIL <= '1';
              FAIL_NUM <= "01110011";
              state <= "11111101";
            ELSE
              state <= "10000001";
            END IF;
            uut_rst <= '0';
          WHEN "10000001" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000110000";
            uut_y <= "000000001010";
            uut_fx <= "1001001000";
            uut_fy <= "0110110001";
            uut_ft <= "0100110100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000010110110010000" OR uut_a_0_1 /= "111101100000111000110010000" OR uut_a_0_2 /= "111100111011100000110000000" OR uut_a_0_3 /= "000000000000001101100000000" OR uut_a_0_4 /= "111110100001101101100000000" OR uut_a_0_5 /= "111110001011100100000000000" OR uut_a_1_0 /= "111111111111110110000011100" OR uut_a_1_1 /= "000001000101011101001101101" OR uut_a_1_2 /= "000001010101110001011001000" OR uut_a_1_3 /= "111111111111111010000110110" OR uut_a_1_4 /= "000000101001001010001100110" OR uut_a_1_5 /= "000000110010110100111110010" OR uut_a_2_0 /= "111111111111110011101110000" OR uut_a_2_1 /= "000001010101110001011001000" OR uut_a_2_2 /= "000001101001111010110110001" OR uut_a_2_3 /= "111111111111111000101110010" OR uut_a_2_4 /= "000000110010110100111110010" OR uut_a_2_5 /= "000000111110110001000110000" OR uut_a_3_0 /= "000000000000001101100000000" OR uut_a_3_1 /= "111110100001101101100000000" OR uut_a_3_2 /= "111110001011100100000000000" OR uut_a_3_3 /= "000000000000001000000000000" OR uut_a_3_4 /= "111111001000001000000000000" OR uut_a_3_5 /= "111110111011000000000000000" OR uut_a_4_0 /= "111111111111111010000110110" OR uut_a_4_1 /= "000000101001001010001100110" OR uut_a_4_2 /= "000000110010110100111110010" OR uut_a_4_3 /= "111111111111111100100000100" OR uut_a_4_4 /= "000000011000011001000000100" OR uut_a_4_5 /= "000000011110000111101100000" OR uut_a_5_0 /= "111111111111111000101110010" OR uut_a_5_1 /= "000000110010110100111110010" OR uut_a_5_2 /= "000000111110110001000110000" OR uut_a_5_3 /= "111111111111111011101100000" OR uut_a_5_4 /= "000000011110000111101100000" OR uut_a_5_5 /= "000000100101001100100000000" THEN
              FAIL <= '1';
              FAIL_NUM <= "01110100";
              state <= "11111101";
            ELSE
              state <= "10000010";
            END IF;
            uut_rst <= '0';
          WHEN "10000010" =>
            uut_coord_shift <= "0101";
            uut_x <= "111111100101";
            uut_y <= "000000000101";
            uut_fx <= "0111110000";
            uut_fy <= "0011011101";
            uut_ft <= "0101011011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000001011101110110" OR uut_a_0_1 /= "000000111100001101100111101" OR uut_a_0_2 /= "111101010110001011010001001" OR uut_a_0_3 /= "000000000000000011110010001" OR uut_a_0_4 /= "000000010011011011000110100" OR uut_a_0_5 /= "111111001001001101111101010" OR uut_a_1_0 /= "000000000000000011110000110" OR uut_a_1_1 /= "000000010011010100001111100" OR uut_a_1_2 /= "111111001001100001010011010" OR uut_a_1_3 /= "000000000000000001001101101" OR uut_a_1_4 /= "000000000110001110110010011" OR uut_a_1_5 /= "111111101110011011010000100" OR uut_a_2_0 /= "111111111111110101011000101" OR uut_a_2_1 /= "111111001001100001010011010" OR uut_a_2_2 /= "000010011001101001110111011" OR uut_a_2_3 /= "111111111111111100100100110" OR uut_a_2_4 /= "111111101110011011010000100" OR uut_a_2_5 /= "000000110001100100001101110" OR uut_a_3_0 /= "000000000000000011110010001" OR uut_a_3_1 /= "000000010011011011000110100" OR uut_a_3_2 /= "111111001001001101111101010" OR uut_a_3_3 /= "000000000000000001001110001" OR uut_a_3_4 /= "000000000110010001000000000" OR uut_a_3_5 /= "111111101110010101000001001" OR uut_a_4_0 /= "000000000000000001001101101" OR uut_a_4_1 /= "000000000110001110110010011" OR uut_a_4_2 /= "111111101110011011010000100" OR uut_a_4_3 /= "000000000000000000011001000" OR uut_a_4_4 /= "000000000010000000101001000" OR uut_a_4_5 /= "111111111010010101001011100" OR uut_a_5_0 /= "111111111111111100100100110" OR uut_a_5_1 /= "111111101110011011010000100" OR uut_a_5_2 /= "000000110001100100001101110" OR uut_a_5_3 /= "111111111111111110111001010" OR uut_a_5_4 /= "111111111010010101001011100" OR uut_a_5_5 /= "000000001111111111010010111" THEN
              FAIL <= '1';
              FAIL_NUM <= "01110101";
              state <= "11111101";
            ELSE
              state <= "10000011";
            END IF;
            uut_rst <= '0';
          WHEN "10000011" =>
            uut_coord_shift <= "0101";
            uut_x <= "111111111000";
            uut_y <= "111111111101";
            uut_fx <= "0000111110";
            uut_fy <= "1100010100";
            uut_ft <= "0011111111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000011000100000000" OR uut_a_0_1 /= "000010101000011100000000000" OR uut_a_0_2 /= "000100010111000100100000000" OR uut_a_0_3 /= "111111111111100110000101000" OR uut_a_0_4 /= "111101001101110010011000000" OR uut_a_0_5 /= "111011011000101110111101000" OR uut_a_1_0 /= "000000000000001010100001110" OR uut_a_1_1 /= "000001001000011000000010000" OR uut_a_1_2 /= "000001110111111010011011110" OR uut_a_1_3 /= "111111111111110100110111001" OR uut_a_1_4 /= "111110110011011011001001010" OR uut_a_1_5 /= "111110000001001000001011001" OR uut_a_2_0 /= "000000000000010001011100010" OR uut_a_2_1 /= "000001110111111010011011110" OR uut_a_2_2 /= "000011000110101011001001000" OR uut_a_2_3 /= "111111111111101101100010111" OR uut_a_2_4 /= "111110000001001000001011001" OR uut_a_2_5 /= "111100101101110010111011010" OR uut_a_3_0 /= "111111111111100110000101000" OR uut_a_3_1 /= "111101001101110010011000000" OR uut_a_3_2 /= "111011011000101110111101000" OR uut_a_3_3 /= "000000000000011011011011010" OR uut_a_3_4 /= "000010111100100011100011110" OR uut_a_3_5 /= "000100111000011001110000000" OR uut_a_4_0 /= "111111111111110100110111001" OR uut_a_4_1 /= "111110110011011011001001010" OR uut_a_4_2 /= "111110000001001000001011001" OR uut_a_4_3 /= "000000000000001011110010001" OR uut_a_4_4 /= "000001010001000001010001110" OR uut_a_4_5 /= "000010000110001111000100001" OR uut_a_5_0 /= "111111111111101101100010111" OR uut_a_5_1 /= "111110000001001000001011001" OR uut_a_5_2 /= "111100101101110010111011010" OR uut_a_5_3 /= "000000000000010011100001100" OR uut_a_5_4 /= "000010000110001111000100001" OR uut_a_5_5 /= "000011011110011001110101010" THEN
              FAIL <= '1';
              FAIL_NUM <= "01110110";
              state <= "11111101";
            ELSE
              state <= "10000100";
            END IF;
            uut_rst <= '0';
          WHEN "10000100" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000000000";
            uut_y <= "000000010010";
            uut_fx <= "1100111011";
            uut_fy <= "1010001110";
            uut_ft <= "1111100111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000011111101001" OR uut_a_0_1 /= "000000101010100111000001101" OR uut_a_0_2 /= "111111010010010001001111100" OR uut_a_0_3 /= "111111111111111001111110101" OR uut_a_0_4 /= "111110111111001000110111000" OR uut_a_0_5 /= "000001000101100111001011010" OR uut_a_1_0 /= "000000000000000010101010011" OR uut_a_1_1 /= "000000011100101100001101110" OR uut_a_1_2 /= "111111100001001101010011000" OR uut_a_1_3 /= "111111111111111011111100100" OR uut_a_1_4 /= "111111010100010100110111110" OR uut_a_1_5 /= "000000101110110111110110001" OR uut_a_2_0 /= "111111111111111101001001000" OR uut_a_2_1 /= "111111100001001101010011000" OR uut_a_2_2 /= "000000100001000011000010100" OR uut_a_2_3 /= "000000000000000100010110011" OR uut_a_2_4 /= "000000101110110111110110001" OR uut_a_2_5 /= "111111001101101100011100000" OR uut_a_3_0 /= "111111111111111001111110101" OR uut_a_3_1 /= "111110111111001000110111000" OR uut_a_3_2 /= "000001000101100111001011010" OR uut_a_3_3 /= "000000000000001001001010100" OR uut_a_3_4 /= "000001100010101110111101010" OR uut_a_3_5 /= "111110010110000010001110111" OR uut_a_4_0 /= "111111111111111011111100100" OR uut_a_4_1 /= "111111010100010100110111110" OR uut_a_4_2 /= "000000101110110111110110001" OR uut_a_4_3 /= "000000000000000110001010111" OR uut_a_4_4 /= "000001000010011110110011100" OR uut_a_4_5 /= "111110111000101001100100001" OR uut_a_5_0 /= "000000000000000100010110011" OR uut_a_5_1 /= "000000101110110111110110001" OR uut_a_5_2 /= "111111001101101100011100000" OR uut_a_5_3 /= "111111111111111001011000001" OR uut_a_5_4 /= "111110111000101001100100001" OR uut_a_5_5 /= "000001001100100100111000110" THEN
              FAIL <= '1';
              FAIL_NUM <= "01110111";
              state <= "11111101";
            ELSE
              state <= "10000101";
            END IF;
            uut_rst <= '0';
          WHEN "10000101" =>
            uut_coord_shift <= "0101";
            uut_x <= "111111101111";
            uut_y <= "000000100100";
            uut_fx <= "0100011111";
            uut_fy <= "0010101101";
            uut_ft <= "1010001001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000100100011000000100000" OR uut_a_0_1 /= "000000000000000000000000000" OR uut_a_0_2 /= "111111101101110011111110000" OR uut_a_0_3 /= "111111110001110111010100000" OR uut_a_0_4 /= "000000000000000000000000000" OR uut_a_0_5 /= "000000000111000100010110000" OR uut_a_1_0 /= "000000000000000000000000000" OR uut_a_1_1 /= "000000000000000000000000000" OR uut_a_1_2 /= "000000000000000000000000000" OR uut_a_1_3 /= "000000000000000000000000000" OR uut_a_1_4 /= "000000000000000000000000000" OR uut_a_1_5 /= "000000000000000000000000000" OR uut_a_2_0 /= "111111111111011011100111111" OR uut_a_2_1 /= "000000000000000000000000000" OR uut_a_2_2 /= "000000000000010010001100000" OR uut_a_2_3 /= "000000000000001110001000101" OR uut_a_2_4 /= "000000000000000000000000000" OR uut_a_2_5 /= "111111111111111000111011101" OR uut_a_3_0 /= "111111110001110111010100000" OR uut_a_3_1 /= "000000000000000000000000000" OR uut_a_3_2 /= "000000000111000100010110000" OR uut_a_3_3 /= "000000000101011111100100000" OR uut_a_3_4 /= "000000000000000000000000000" OR uut_a_3_5 /= "111111111101010000001110000" OR uut_a_4_0 /= "000000000000000000000000000" OR uut_a_4_1 /= "000000000000000000000000000" OR uut_a_4_2 /= "000000000000000000000000000" OR uut_a_4_3 /= "000000000000000000000000000" OR uut_a_4_4 /= "000000000000000000000000000" OR uut_a_4_5 /= "000000000000000000000000000" OR uut_a_5_0 /= "000000000000001110001000101" OR uut_a_5_1 /= "000000000000000000000000000" OR uut_a_5_2 /= "111111111111111000111011101" OR uut_a_5_3 /= "111111111111111010100000011" OR uut_a_5_4 /= "000000000000000000000000000" OR uut_a_5_5 /= "000000000000000010101111110" THEN
              FAIL <= '1';
              FAIL_NUM <= "01111000";
              state <= "11111101";
            ELSE
              state <= "10000110";
            END IF;
            uut_rst <= '0';
          WHEN "10000110" =>
            uut_coord_shift <= "0101";
            uut_x <= "111111000011";
            uut_y <= "000000000111";
            uut_fx <= "1100110100";
            uut_fy <= "0111000010";
            uut_ft <= "0111101100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000111001001100010000000" OR uut_a_0_1 /= "011010010111001001011000000" OR uut_a_0_2 /= "100110000101011100110000000" OR uut_a_0_3 /= "111111011010011011001000000" OR uut_a_0_4 /= "101110101011100000001100000" OR uut_a_0_5 /= "010001000001101101011000000" OR uut_a_1_0 /= "000000110100101110010010110" OR uut_a_1_1 /= "011000010011010101101001001" OR uut_a_1_2 /= "101000000111000001100000010" OR uut_a_1_3 /= "111111011101010111000000011" OR uut_a_1_4 /= "110000000010000110101011000" OR uut_a_1_5 /= "001111101100100100110101001" OR uut_a_2_0 /= "111111001100001010111001100" OR uut_a_2_1 /= "101000000111000001100000010" OR uut_a_2_2 /= "010111011111000011111100100" OR uut_a_2_3 /= "000000100010000011011010110" OR uut_a_2_4 /= "001111101100100100110101001" OR uut_a_2_5 /= "110000100100011100111000010" OR uut_a_3_0 /= "111111011010011011001000000" OR uut_a_3_1 /= "101110101011100000001100000" OR uut_a_3_2 /= "010001000001101101011000000" OR uut_a_3_3 /= "000000011000101100000100000" OR uut_a_3_4 /= "001011011000010011110110000" OR uut_a_3_5 /= "110100110100000010001100000" OR uut_a_4_0 /= "111111011101010111000000011" OR uut_a_4_1 /= "110000000010000110101011000" OR uut_a_4_2 /= "001111101100100100110101001" OR uut_a_4_3 /= "000000010110110000100111101" OR uut_a_4_4 /= "001010011111011010010010110" OR uut_a_4_5 /= "110101101011111110000001000" OR uut_a_5_0 /= "000000100010000011011010110" OR uut_a_5_1 /= "001111101100100100110101001" OR uut_a_5_2 /= "110000100100011100111000010" OR uut_a_5_3 /= "111111101001101000000100011" OR uut_a_5_4 /= "110101101011111110000001000" OR uut_a_5_5 /= "001010001000110110000001001" THEN
              FAIL <= '1';
              FAIL_NUM <= "01111001";
              state <= "11111101";
            ELSE
              state <= "10000111";
            END IF;
            uut_rst <= '0';
          WHEN "10000111" =>
            uut_coord_shift <= "0101";
            uut_x <= "111111100101";
            uut_y <= "000000100110";
            uut_fx <= "0110010110";
            uut_fy <= "0001100100";
            uut_ft <= "0110001001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000100111011000100000" OR uut_a_0_1 /= "000000011011000100110110000" OR uut_a_0_2 /= "000000110110001001101100000" OR uut_a_0_3 /= "111111111011101111000110000" OR uut_a_0_4 /= "111111101000100011000001000" OR uut_a_0_5 /= "111111010001000110000010000" OR uut_a_1_0 /= "000000000000110110001001101" OR uut_a_1_1 /= "000000000100101001110101010" OR uut_a_1_2 /= "000000001001010011101010100" OR uut_a_1_3 /= "111111111111010001000110000" OR uut_a_1_4 /= "111111111011111110000001001" OR uut_a_1_5 /= "111111110111111100000010010" OR uut_a_2_0 /= "000000000001101100010011011" OR uut_a_2_1 /= "000000001001010011101010100" OR uut_a_2_2 /= "000000010010100111010101001" OR uut_a_2_3 /= "111111111110100010001100000" OR uut_a_2_4 /= "111111110111111100000010010" OR uut_a_2_5 /= "111111101111111000000100101" OR uut_a_3_0 /= "111111111011101111000110000" OR uut_a_3_1 /= "111111101000100011000001000" OR uut_a_3_2 /= "111111010001000110000010000" OR uut_a_3_3 /= "000000000011101100011001000" OR uut_a_3_4 /= "000000010100010100001001100" OR uut_a_3_5 /= "000000101000101000010011000" OR uut_a_4_0 /= "111111111111010001000110000" OR uut_a_4_1 /= "111111111011111110000001001" OR uut_a_4_2 /= "111111110111111100000010010" OR uut_a_4_3 /= "000000000000101000101000010" OR uut_a_4_4 /= "000000000011011111011101101" OR uut_a_4_5 /= "000000000110111110111011010" OR uut_a_5_0 /= "111111111110100010001100000" OR uut_a_5_1 /= "111111110111111100000010010" OR uut_a_5_2 /= "111111101111111000000100101" OR uut_a_5_3 /= "000000000001010001010000100" OR uut_a_5_4 /= "000000000110111110111011010" OR uut_a_5_5 /= "000000001101111101110110100" THEN
              FAIL <= '1';
              FAIL_NUM <= "01111010";
              state <= "11111101";
            ELSE
              state <= "10001000";
            END IF;
            uut_rst <= '0';
          WHEN "10001000" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000111000";
            uut_y <= "000000000110";
            uut_fx <= "0011101010";
            uut_fy <= "0001001111";
            uut_ft <= "1000011010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000111001101010100100000" OR uut_a_0_1 /= "100100100001001101110110000" OR uut_a_0_2 /= "101000000111111000000110000" OR uut_a_0_3 /= "000000010010011001000010000" OR uut_a_0_4 /= "110111001111000100100011000" OR uut_a_0_5 /= "111000011000101000101011000" OR uut_a_1_0 /= "111111001001000010011011101" OR uut_a_1_1 /= "011010001100010101110011100" OR uut_a_1_2 /= "010110110000011111100010010" OR uut_a_1_3 /= "111111101110011110001001000" OR uut_a_1_4 /= "001000010110101000101010101" OR uut_a_1_5 /= "000111010000100001001111000" OR uut_a_2_0 /= "111111010000001111110000001" OR uut_a_2_1 /= "010110110000011111100010010" OR uut_a_2_2 /= "010011110001011110100011000" OR uut_a_2_3 /= "111111110000110001010001010" OR uut_a_2_4 /= "000111010000100001001111000" OR uut_a_2_5 /= "000110010011100110010100011" OR uut_a_3_0 /= "000000010010011001000010000" OR uut_a_3_1 /= "110111001111000100100011000" OR uut_a_3_2 /= "111000011000101000101011000" OR uut_a_3_3 /= "000000000101110111011001000" OR uut_a_3_4 /= "111101001101000110100101100" OR uut_a_3_5 /= "111101100100100100001001100" OR uut_a_4_0 /= "111111101110011110001001000" OR uut_a_4_1 /= "001000010110101000101010101" OR uut_a_4_2 /= "000111010000100001001111000" OR uut_a_4_3 /= "111111111010011010001101001" OR uut_a_4_4 /= "000010101010100000101110010" OR uut_a_4_5 /= "000010010100001001100010111" OR uut_a_5_0 /= "111111110000110001010001010" OR uut_a_5_1 /= "000111010000100001001111000" OR uut_a_5_2 /= "000110010011100110010100011" OR uut_a_5_3 /= "111111111011001001001000010" OR uut_a_5_4 /= "000010010100001001100010111" OR uut_a_5_5 /= "000010000000101110000100001" THEN
              FAIL <= '1';
              FAIL_NUM <= "01111011";
              state <= "11111101";
            ELSE
              state <= "10001001";
            END IF;
            uut_rst <= '0';
          WHEN "10001001" =>
            uut_coord_shift <= "0101";
            uut_x <= "111111111010";
            uut_y <= "000000010010";
            uut_fx <= "0000010110";
            uut_fy <= "1101111101";
            uut_ft <= "0111000000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000001101101101101001000" OR uut_a_0_1 /= "111110101101101110001010000" OR uut_a_0_2 /= "111010110110111000101000000" OR uut_a_0_3 /= "000000001110010110011000000" OR uut_a_0_4 /= "111110101001111001110000000" OR uut_a_0_5 /= "111010100111100111000000000" OR uut_a_1_0 /= "111111111101011011011100010" OR uut_a_1_1 /= "000000001111011011010110001" OR uut_a_1_2 /= "000000111101101101011000100" OR uut_a_1_3 /= "111111111101010011110011100" OR uut_a_1_4 /= "000000010000001001001011000" OR uut_a_1_5 /= "000001000000100100101100000" OR uut_a_2_0 /= "111111110101101101110001010" OR uut_a_2_1 /= "000000111101101101011000100" OR uut_a_2_2 /= "000011110110110101100010000" OR uut_a_2_3 /= "111111110101001111001110000" OR uut_a_2_4 /= "000001000000100100101100000" OR uut_a_2_5 /= "000100000010010010110000000" OR uut_a_3_0 /= "000000001110010110011000000" OR uut_a_3_1 /= "111110101001111001110000000" OR uut_a_3_2 /= "111010100111100111000000000" OR uut_a_3_3 /= "000000001111000001000000000" OR uut_a_3_4 /= "111110100101111010000000000" OR uut_a_3_5 /= "111010010111101000000000000" OR uut_a_4_0 /= "111111111101010011110011100" OR uut_a_4_1 /= "000000010000001001001011000" OR uut_a_4_2 /= "000001000000100100101100000" OR uut_a_4_3 /= "111111111101001011110100000" OR uut_a_4_4 /= "000000010000111001001000000" OR uut_a_4_5 /= "000001000011100100100000000" OR uut_a_5_0 /= "111111110101001111001110000" OR uut_a_5_1 /= "000001000000100100101100000" OR uut_a_5_2 /= "000100000010010010110000000" OR uut_a_5_3 /= "111111110100101111010000000" OR uut_a_5_4 /= "000001000011100100100000000" OR uut_a_5_5 /= "000100001110010010000000000" THEN
              FAIL <= '1';
              FAIL_NUM <= "01111100";
              state <= "11111101";
            ELSE
              state <= "10001010";
            END IF;
            uut_rst <= '0';
          WHEN "10001010" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000101010";
            uut_y <= "000000101100";
            uut_fx <= "1101111101";
            uut_fy <= "0001011111";
            uut_ft <= "0101111101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000100100100100001001000" OR uut_a_0_1 /= "110011011011100100111010000" OR uut_a_0_2 /= "111010100100101000101010100" OR uut_a_0_3 /= "111111011010110111100101000" OR uut_a_0_4 /= "001100110000111001010010000" OR uut_a_0_5 /= "000101100000110000000000100" OR uut_a_1_0 /= "111111100110110111001001110" OR uut_a_1_1 /= "001000101001000010101000001" OR uut_a_1_2 /= "000011101110110100000010110" OR uut_a_1_3 /= "000000011001100001110010100" OR uut_a_1_4 /= "110111001110011000100111101" OR uut_a_1_5 /= "111100001101011110111111101" OR uut_a_2_0 /= "111111110101001001010001010" OR uut_a_2_1 /= "000011101110110100000010110" OR uut_a_2_2 /= "000001100111000111111011011" OR uut_a_2_3 /= "000000001011000001100000000" OR uut_a_2_4 /= "111100001101011110111111101" OR uut_a_2_5 /= "111110010111010001101111110" OR uut_a_3_0 /= "111111011010110111100101000" OR uut_a_3_1 /= "001100110000111001010010000" OR uut_a_3_2 /= "000101100000110000000000100" OR uut_a_3_3 /= "000000100101101101010001000" OR uut_a_3_4 /= "110011000010011100001010000" OR uut_a_3_5 /= "111010011001110001111110100" OR uut_a_4_0 /= "000000011001100001110010100" OR uut_a_4_1 /= "110111001110011000100111101" OR uut_a_4_2 /= "111100001101011110111111101" OR uut_a_4_3 /= "111111100110000100111000010" OR uut_a_4_4 /= "001000111010010100101001001" OR uut_a_4_5 /= "000011110110010001101001000" OR uut_a_5_0 /= "000000001011000001100000000" OR uut_a_5_1 /= "111100001101011110111111101" OR uut_a_5_2 /= "111110010111010001101111110" OR uut_a_5_3 /= "111111110100110011100011111" OR uut_a_5_4 /= "000011110110010001101001000" OR uut_a_5_5 /= "000001101010010110001010011" THEN
              FAIL <= '1';
              FAIL_NUM <= "01111101";
              state <= "11111101";
            ELSE
              state <= "10001011";
            END IF;
            uut_rst <= '0';
          WHEN "10001011" =>
            uut_coord_shift <= "0101";
            uut_x <= "000000110111";
            uut_y <= "000000010101";
            uut_fx <= "1011010100";
            uut_fy <= "0010011110";
            uut_ft <= "1001001010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000110100010101100001000" OR uut_a_0_1 /= "010110011111001111101011100" OR uut_a_0_2 /= "111011000101111110111010000" OR uut_a_0_3 /= "000000010010001100101111000" OR uut_a_0_4 /= "000111110100011110001100100" OR uut_a_0_5 /= "111110010010110011100110000" OR uut_a_1_0 /= "000000101100111110011111010" OR uut_a_1_1 /= "010011010100110110011110011" OR uut_a_1_2 /= "111011110010001001000011110" OR uut_a_1_3 /= "000000001111101000111100011" OR uut_a_1_4 /= "000110101110000101111100101" OR uut_a_1_5 /= "111110100010001010010101101" OR uut_a_2_0 /= "111111110110001011111101110" OR uut_a_2_1 /= "111011110010001001000011110" OR uut_a_2_2 /= "000000111010111000001101001" OR uut_a_2_3 /= "111111111100100101100111001" OR uut_a_2_4 /= "111110100010001010010101101" OR uut_a_2_5 /= "000000010100011110010100111" OR uut_a_3_0 /= "000000010010001100101111000" OR uut_a_3_1 /= "000111110100011110001100100" OR uut_a_3_2 /= "111110010010110011100110000" OR uut_a_3_3 /= "000000000110010101000001000" OR uut_a_3_4 /= "000010101110000001111011100" OR uut_a_3_5 /= "111111011010000001111010000" OR uut_a_4_0 /= "000000001111101000111100011" OR uut_a_4_1 /= "000110101110000101111100101" OR uut_a_4_2 /= "111110100010001010010101101" OR uut_a_4_3 /= "000000000101011100000011110" OR uut_a_4_4 /= "000010010101100011101010001" OR uut_a_4_5 /= "111111011111010111101000110" OR uut_a_5_0 /= "111111111100100101100111001" OR uut_a_5_1 /= "111110100010001010010101101" OR uut_a_5_2 /= "000000010100011110010100111" OR uut_a_5_3 /= "111111111110110100000011110" OR uut_a_5_4 /= "111111011111010111101000110" OR uut_a_5_5 /= "000000000111000111101001001" THEN
              FAIL <= '1';
              FAIL_NUM <= "01111110";
              state <= "11111101";
            ELSE
              state <= "10001100";
            END IF;
            uut_rst <= '0';
          WHEN "10001100" =>
            uut_coord_shift <= "0110";
            uut_x <= "111111101001";
            uut_y <= "000000101010";
            uut_fx <= "0110111100";
            uut_fy <= "0100111110";
            uut_ft <= "1111110000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000001000111010000001000" OR uut_a_0_1 /= "000010100100110001010010100" OR uut_a_0_2 /= "000000010110010001000010100" OR uut_a_0_3 /= "000000010010110010101101000" OR uut_a_0_4 /= "000101011011101010000000100" OR uut_a_0_5 /= "000000101110111110110000100" OR uut_a_1_0 /= "000000000101001001100010100" OR uut_a_1_1 /= "000001011111010000011111101" OR uut_a_1_2 /= "000000001100110111110110011" OR uut_a_1_3 /= "000000001010110111010100000" OR uut_a_1_4 /= "000011001000111111010010010" OR uut_a_1_5 /= "000000011011001010010010000" OR uut_a_2_0 /= "000000000000101100100010000" OR uut_a_2_1 /= "000000001100110111110110011" OR uut_a_2_2 /= "000000000001101111010101001" OR uut_a_2_3 /= "000000000001011101111101100" OR uut_a_2_4 /= "000000011011001010010010000" OR uut_a_2_5 /= "000000000011101010111001110" OR uut_a_3_0 /= "000000010010110010101101000" OR uut_a_3_1 /= "000101011011101010000000100" OR uut_a_3_2 /= "000000101110111110110000100" OR uut_a_3_3 /= "000000100111101001101001000" OR uut_a_3_4 /= "001011011101100010010110100" OR uut_a_3_5 /= "000001100011001000000110100" OR uut_a_4_0 /= "000000001010110111010100000" OR uut_a_4_1 /= "000011001000111111010010010" OR uut_a_4_2 /= "000000011011001010010010000" OR uut_a_4_3 /= "000000010110111011000100101" OR uut_a_4_4 /= "000110101000000100110111000" OR uut_a_4_5 /= "000000111001010011101011110" OR uut_a_5_0 /= "000000000001011101111101100" OR uut_a_5_1 /= "000000011011001010010010000" OR uut_a_5_2 /= "000000000011101010111001110" OR uut_a_5_3 /= "000000000011000110010000001" OR uut_a_5_4 /= "000000111001010011101011110" OR uut_a_5_5 /= "000000000111101111101000100" THEN
              FAIL <= '1';
              FAIL_NUM <= "01111111";
              state <= "11111101";
            ELSE
              state <= "10001101";
            END IF;
            uut_rst <= '0';
          WHEN "10001101" =>
            uut_coord_shift <= "0110";
            uut_x <= "000001000001";
            uut_y <= "111111101011";
            uut_fx <= "0111100011";
            uut_fy <= "0111110100";
            uut_ft <= "0101110101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000010111110001000000000" OR uut_a_0_1 /= "111011010110111011100000000" OR uut_a_0_2 /= "110101001110110011000000000" OR uut_a_0_3 /= "111111101110110111001000000" OR uut_a_0_4 /= "000011010110001110111100000" OR uut_a_0_5 /= "000111110001000001011000000" OR uut_a_1_0 /= "111111110110101101110111000" OR uut_a_1_1 /= "000001110100000010110000100" OR uut_a_1_2 /= "000100001101001110000101000" OR uut_a_1_3 /= "000000000110101100011101111" OR uut_a_1_4 /= "111110101100010100001010100" OR uut_a_1_5 /= "111100111101110110011101101" OR uut_a_2_0 /= "111111101010011101100110000" OR uut_a_2_1 /= "000100001101001110000101000" OR uut_a_2_2 /= "001001110000100101110010000" OR uut_a_2_3 /= "000000001111100010000010110" OR uut_a_2_4 /= "111100111101110110011101101" OR uut_a_2_5 /= "111000111101100100110000010" OR uut_a_3_0 /= "111111101110110111001000000" OR uut_a_3_1 /= "000011010110001110111100000" OR uut_a_3_2 /= "000111110001000001011000000" OR uut_a_3_3 /= "000000001100010111000001000" OR uut_a_3_4 /= "111101100101100000010011100" OR uut_a_3_5 /= "111010011001100100100011000" OR uut_a_4_0 /= "000000000110101100011101111" OR uut_a_4_1 /= "111110101100010100001010100" OR uut_a_4_2 /= "111100111101110110011101101" OR uut_a_4_3 /= "111111111011001011000000100" OR uut_a_4_4 /= "000000111100010110011000011" OR uut_a_4_5 /= "000010001100000000101110010" OR uut_a_5_0 /= "000000001111100010000010110" OR uut_a_5_1 /= "111100111101110110011101101" OR uut_a_5_2 /= "111000111101100100110000010" OR uut_a_5_3 /= "111111110100110011001001000" OR uut_a_5_4 /= "000010001100000000101110010" OR uut_a_5_5 /= "000101000100110100111000010" THEN
              FAIL <= '1';
              FAIL_NUM <= "10000000";
              state <= "11111101";
            ELSE
              state <= "10001110";
            END IF;
            uut_rst <= '0';
          WHEN "10001110" =>
            uut_coord_shift <= "0110";
            uut_x <= "111111100100";
            uut_y <= "111111110101";
            uut_fx <= "1011111101";
            uut_fy <= "0100100011";
            uut_ft <= "0110001000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000101111010001000000000" OR uut_a_0_1 /= "010001101110011000000000000" OR uut_a_0_2 /= "000011101100010101000000000" OR uut_a_0_3 /= "111111010001011111001000000" OR uut_a_0_4 /= "101110100011101011000000000" OR uut_a_0_5 /= "111100010111011011101000000" OR uut_a_1_0 /= "000000100011011100110000000" OR uut_a_1_1 /= "001101010010110010000000000" OR uut_a_1_2 /= "000010110001001111110000000" OR uut_a_1_3 /= "111111011101000111010110000" OR uut_a_1_4 /= "110010111010110000010000000" OR uut_a_1_5 /= "111101010001100100101110000" OR uut_a_2_0 /= "000000000111011000101010000" OR uut_a_2_1 /= "000010110001001111110000000" OR uut_a_2_2 /= "000000100100111011010010000" OR uut_a_2_3 /= "111111111000101110110111010" OR uut_a_2_4 /= "111101010001100100101110000" OR uut_a_2_5 /= "111111011011101010010100010" OR uut_a_3_0 /= "111111010001011111001000000" OR uut_a_3_1 /= "101110100011101011000000000" OR uut_a_3_2 /= "111100010111011011101000000" OR uut_a_3_3 /= "000000101101110001100001000" OR uut_a_3_4 /= "010001001010100100011000000" OR uut_a_3_5 /= "000011100100110111100101000" OR uut_a_4_0 /= "111111011101000111010110000" OR uut_a_4_1 /= "110010111010110000010000000" OR uut_a_4_2 /= "111101010001100100101110000" OR uut_a_4_3 /= "000000100010010101001000110" OR uut_a_4_4 /= "001100110111111011010010000" OR uut_a_4_5 /= "000010101011101001101011110" OR uut_a_5_0 /= "111111111000101110110111010" OR uut_a_5_1 /= "111101010001100100101110000" OR uut_a_5_2 /= "111111011011101010010100010" OR uut_a_5_3 /= "000000000111001001101111001" OR uut_a_5_4 /= "000010101011101001101011110" OR uut_a_5_5 /= "000000100011110000101011110" THEN
              FAIL <= '1';
              FAIL_NUM <= "10000001";
              state <= "11111101";
            ELSE
              state <= "10001111";
            END IF;
            uut_rst <= '0';
          WHEN "10001111" =>
            uut_coord_shift <= "0110";
            uut_x <= "000001101001";
            uut_y <= "000000001110";
            uut_fx <= "0001100101";
            uut_fy <= "1010011000";
            uut_ft <= "0110011001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000111100000100000000000" OR uut_a_0_1 /= "110011010101001010000000000" OR uut_a_0_2 /= "000010010110001010000000000" OR uut_a_0_3 /= "000000011010110000110000000" OR uut_a_0_4 /= "111010010110101101111000000" OR uut_a_0_5 /= "000001000010111001111000000" OR uut_a_1_0 /= "111111100110101010010100000" OR uut_a_1_1 /= "000101010110000100110010000" OR uut_a_1_2 /= "111111000000101001110010000" OR uut_a_1_3 /= "111111110100101101011011110" OR uut_a_1_4 /= "000010011000011010101001011" OR uut_a_1_5 /= "111111100011110001100101011" OR uut_a_2_0 /= "000000000100101100010100000" OR uut_a_2_1 /= "111111000000101001110010000" OR uut_a_2_2 /= "000000001011101110110010000" OR uut_a_2_3 /= "000000000010000101110011110" OR uut_a_2_4 /= "111111100011110001100101011" OR uut_a_2_5 /= "000000000101001110100001011" OR uut_a_3_0 /= "000000011010110000110000000" OR uut_a_3_1 /= "111010010110101101111000000" OR uut_a_3_2 /= "000001000010111001111000000" OR uut_a_3_3 /= "000000001011111011001001000" OR uut_a_3_4 /= "111101011111000001100110100" OR uut_a_3_5 /= "000000011101110011110110100" OR uut_a_4_0 /= "111111110100101101011011110" OR uut_a_4_1 /= "000010011000011010101001011" OR uut_a_4_2 /= "111111100011110001100101011" OR uut_a_4_3 /= "111111111010111110000011001" OR uut_a_4_4 /= "000001000011111010010100110" OR uut_a_4_5 /= "111111110011011011001000000" OR uut_a_5_0 /= "000000000010000101110011110" OR uut_a_5_1 /= "111111100011110001100101011" OR uut_a_5_2 /= "000000000101001110100001011" OR uut_a_5_3 /= "000000000000111011100111101" OR uut_a_5_4 /= "111111110011011011001000000" OR uut_a_5_5 /= "000000000010010101000011010" THEN
              FAIL <= '1';
              FAIL_NUM <= "10000010";
              state <= "11111101";
            ELSE
              state <= "10010000";
            END IF;
            uut_rst <= '0';
          WHEN "10010000" =>
            uut_coord_shift <= "0110";
            uut_x <= "111111110100";
            uut_y <= "111110110101";
            uut_fx <= "0110011001";
            uut_fy <= "0100001101";
            uut_ft <= "0110001000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000111100000100000" OR uut_a_0_1 /= "111111111100001111110000000" OR uut_a_0_2 /= "111111111110100101111010000" OR uut_a_0_3 /= "111111111100011011011000000" OR uut_a_0_4 /= "000000001110010010100000000" OR uut_a_0_5 /= "000000000101010110111100000" OR uut_a_1_0 /= "111111111111111000011111100" OR uut_a_1_1 /= "000000000000011110000010000" OR uut_a_1_2 /= "000000000000001011010000110" OR uut_a_1_3 /= "000000000000011100100101000" OR uut_a_1_4 /= "111111111110001101101100000" OR uut_a_1_5 /= "111111111111010101001000100" OR uut_a_2_0 /= "111111111111111101001011110" OR uut_a_2_1 /= "000000000000001011010000110" OR uut_a_2_2 /= "000000000000000100001110010" OR uut_a_2_3 /= "000000000000001010101101111" OR uut_a_2_4 /= "111111111111010101001000100" OR uut_a_2_5 /= "111111111111101111111011001" OR uut_a_3_0 /= "111111111100011011011000000" OR uut_a_3_1 /= "000000001110010010100000000" OR uut_a_3_2 /= "000000000101010110111100000" OR uut_a_3_3 /= "000000001101100110010000000" OR uut_a_3_4 /= "111111001001100111000000000" OR uut_a_3_5 /= "111111101011100110101000000" OR uut_a_4_0 /= "000000000000011100100101000" OR uut_a_4_1 /= "111111111110001101101100000" OR uut_a_4_2 /= "111111111111010101001000100" OR uut_a_4_3 /= "111111111110010011001110000" OR uut_a_4_4 /= "000000000110110011001000000" OR uut_a_4_5 /= "000000000010100011001011000" OR uut_a_5_0 /= "000000000000001010101101111" OR uut_a_5_1 /= "111111111111010101001000100" OR uut_a_5_2 /= "111111111111101111111011001" OR uut_a_5_3 /= "111111111111010111001101010" OR uut_a_5_4 /= "000000000010100011001011000" OR uut_a_5_5 /= "000000000000111101001100001" THEN
              FAIL <= '1';
              FAIL_NUM <= "10000011";
              state <= "11111101";
            ELSE
              state <= "10010001";
            END IF;
            uut_rst <= '0';
          WHEN "10010001" =>
            uut_coord_shift <= "0110";
            uut_x <= "111111001001";
            uut_y <= "000000101100";
            uut_fx <= "0010101000";
            uut_fy <= "1001111110";
            uut_ft <= "1110100001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000001001011110011001000" OR uut_a_0_1 /= "000000000000000000000000000" OR uut_a_0_2 /= "000001010101010001100001000" OR uut_a_0_3 /= "000000010001110010111010000" OR uut_a_0_4 /= "000000000000000000000000000" OR uut_a_0_5 /= "000010100000001010001010000" OR uut_a_1_0 /= "000000000000000000000000000" OR uut_a_1_1 /= "000000000000000000000000000" OR uut_a_1_2 /= "000000000000000000000000000" OR uut_a_1_3 /= "000000000000000000000000000" OR uut_a_1_4 /= "000000000000000000000000000" OR uut_a_1_5 /= "000000000000000000000000000" OR uut_a_2_0 /= "000000000010101010100011000" OR uut_a_2_1 /= "000000000000000000000000000" OR uut_a_2_2 /= "000000010111111110111011010" OR uut_a_2_3 /= "000000000101000000010100010" OR uut_a_2_4 /= "000000000000000000000000000" OR uut_a_2_5 /= "000000101101000010110110110" OR uut_a_3_0 /= "000000010001110010111010000" OR uut_a_3_1 /= "000000000000000000000000000" OR uut_a_3_2 /= "000010100000001010001010000" OR uut_a_3_3 /= "000000100001011011000100000" OR uut_a_3_4 /= "000000000000000000000000000" OR uut_a_3_5 /= "000100101100110011100100000" OR uut_a_4_0 /= "000000000000000000000000000" OR uut_a_4_1 /= "000000000000000000000000000" OR uut_a_4_2 /= "000000000000000000000000000" OR uut_a_4_3 /= "000000000000000000000000000" OR uut_a_4_4 /= "000000000000000000000000000" OR uut_a_4_5 /= "000000000000000000000000000" OR uut_a_5_0 /= "000000000101000000010100010" OR uut_a_5_1 /= "000000000000000000000000000" OR uut_a_5_2 /= "000000101101000010110110110" OR uut_a_5_3 /= "000000001001011001100111001" OR uut_a_5_4 /= "000000000000000000000000000" OR uut_a_5_5 /= "000001010100100110100000001" THEN
              FAIL <= '1';
              FAIL_NUM <= "10000100";
              state <= "11111101";
            ELSE
              state <= "10010010";
            END IF;
            uut_rst <= '0';
          WHEN "10010010" =>
            uut_coord_shift <= "0110";
            uut_x <= "111111000111";
            uut_y <= "000000110111";
            uut_fx <= "1100100010";
            uut_fy <= "0110010110";
            uut_ft <= "0101001110";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000010100000111000001000" OR uut_a_0_1 /= "111101010101000100010111100" OR uut_a_0_2 /= "000101101001111110010010000" OR uut_a_0_3 /= "000000001100000111110011000" OR uut_a_0_4 /= "111110011000111101101110100" OR uut_a_0_5 /= "000011011010001100010110000" OR uut_a_1_0 /= "111111111010101010001000101" OR uut_a_1_1 /= "000000101101011001110101110" OR uut_a_1_2 /= "111110011111110110011101001" OR uut_a_1_3 /= "111111111100110001111011011" OR uut_a_1_4 /= "000000011011010111100110101" OR uut_a_1_5 /= "111111000110000010101110001" OR uut_a_2_0 /= "000000001011010011111100100" OR uut_a_2_1 /= "111110011111110110011101001" OR uut_a_2_2 /= "000011001011100111000010001" OR uut_a_2_3 /= "000000000110110100011000101" OR uut_a_2_4 /= "111111000110000010101110001" OR uut_a_2_5 /= "000001111010101110111100011" OR uut_a_3_0 /= "000000001100000111110011000" OR uut_a_3_1 /= "111110011000111101101110100" OR uut_a_3_2 /= "000011011010001100010110000" OR uut_a_3_3 /= "000000000111010011101001000" OR uut_a_3_4 /= "111111000001111001000011100" OR uut_a_3_5 /= "000010000011100001100010000" OR uut_a_4_0 /= "111111111100110001111011011" OR uut_a_4_1 /= "000000011011010111100110101" OR uut_a_4_2 /= "111111000110000010101110001" OR uut_a_4_3 /= "111111111110000011110010000" OR uut_a_4_4 /= "000000010000011111110110000" OR uut_a_4_5 /= "111111011101000100000101111" OR uut_a_5_0 /= "000000000110110100011000101" OR uut_a_5_1 /= "111111000110000010101110001" OR uut_a_5_2 /= "000001111010101110111100011" OR uut_a_5_3 /= "000000000100000111000011000" OR uut_a_5_4 /= "111111011101000100000101111" OR uut_a_5_5 /= "000001001001111110110111001" THEN
              FAIL <= '1';
              FAIL_NUM <= "10000101";
              state <= "11111101";
            ELSE
              state <= "10010011";
            END IF;
            uut_rst <= '0';
          WHEN "10010011" =>
            uut_coord_shift <= "0110";
            uut_x <= "111111100100";
            uut_y <= "000000000000";
            uut_fx <= "0011000111";
            uut_fy <= "0101010110";
            uut_ft <= "0001110000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000001010001010010000000" OR uut_a_0_1 /= "111011001010000111011000000" OR uut_a_0_2 /= "000000100011100011111000000" OR uut_a_0_3 /= "111111101001100101101000000" OR uut_a_0_4 /= "001010101011100100011100000" OR uut_a_0_5 /= "111110110001100011101100000" OR uut_a_1_0 /= "111111110110010100001110110" OR uut_a_1_1 /= "000100100111010110111110001" OR uut_a_1_2 /= "111111011110000110110011101" OR uut_a_1_3 /= "000000010101010111001000111" OR uut_a_1_4 /= "110101110100011110010001010" OR uut_a_1_5 /= "000001001010110000111111000" OR uut_a_2_0 /= "000000000001000111000111110" OR uut_a_2_1 /= "111111011110000110110011101" OR uut_a_2_2 /= "000000000011111000111011001" OR uut_a_2_3 /= "111111111101100011000111011" OR uut_a_2_4 /= "000001001010110000111111000" OR uut_a_2_5 /= "111111110111011010111001110" OR uut_a_3_0 /= "111111101001100101101000000" OR uut_a_3_1 /= "001010101011100100011100000" OR uut_a_3_2 /= "111110110001100011101100000" OR uut_a_3_3 /= "000000110001011100000100000" OR uut_a_3_4 /= "101000011100001000000110000" OR uut_a_3_5 /= "000010101101000010001110000" OR uut_a_4_0 /= "000000010101010111001000111" OR uut_a_4_1 /= "110101110100011110010001010" OR uut_a_4_2 /= "000001001010110000111111000" OR uut_a_4_3 /= "111111010000111000010000001" OR uut_a_4_4 /= "010110011101001100010010010" OR uut_a_4_5 /= "111101011011000100111000101" OR uut_a_5_0 /= "111111111101100011000111011" OR uut_a_5_1 /= "000001001010110000111111000" OR uut_a_5_2 /= "111111110111011010111001110" OR uut_a_5_3 /= "000000000101011010000100011" OR uut_a_5_4 /= "111101011011000100111000101" OR uut_a_5_5 /= "000000010010111011001111100" THEN
              FAIL <= '1';
              FAIL_NUM <= "10000110";
              state <= "11111101";
            ELSE
              state <= "10010100";
            END IF;
            uut_rst <= '0';
          WHEN "10010100" =>
            uut_coord_shift <= "0110";
            uut_x <= "000000010011";
            uut_y <= "111111010100";
            uut_fx <= "1111010011";
            uut_fy <= "0011011011";
            uut_ft <= "0110001010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000101000001111100100000" OR uut_a_0_1 /= "110111100000101101111010000" OR uut_a_0_2 /= "001011111100100111101100000" OR uut_a_0_3 /= "000000001001111010011000000" OR uut_a_0_4 /= "111101111010001011111100000" OR uut_a_0_5 /= "000010111100010101001000000" OR uut_a_1_0 /= "111111101111000001011011110" OR uut_a_1_1 /= "000011100101001100101000100" OR uut_a_1_2 /= "111010111101011011010000011" OR uut_a_1_3 /= "111111111011110100010111111" OR uut_a_1_4 /= "000000111000011100111101101" OR uut_a_1_5 /= "111110110000100011000101101" OR uut_a_2_0 /= "000000010111111001001111011" OR uut_a_2_1 /= "111010111101011011010000011" OR uut_a_2_2 /= "000111000101111111100100001" OR uut_a_2_3 /= "000000000101111000101010010" OR uut_a_2_4 /= "111110110000100011000101101" OR uut_a_2_5 /= "000001101111110100100010110" OR uut_a_3_0 /= "000000001001111010011000000" OR uut_a_3_1 /= "111101111010001011111100000" OR uut_a_3_2 /= "000010111100010101001000000" OR uut_a_3_3 /= "000000000010011100010000000" OR uut_a_3_4 /= "111111011111000010101000000" OR uut_a_3_5 /= "000000101110011000110000000" OR uut_a_4_0 /= "111111111011110100010111111" OR uut_a_4_1 /= "000000111000011100111101101" OR uut_a_4_2 /= "111110110000100011000101101" OR uut_a_4_3 /= "111111111110111110000101010" OR uut_a_4_4 /= "000000001101111001111001001" OR uut_a_4_5 /= "111111101100011011100011110" OR uut_a_5_0 /= "000000000101111000101010010" OR uut_a_5_1 /= "111110110000100011000101101" OR uut_a_5_2 /= "000001101111110100100010110" OR uut_a_5_3 /= "000000000001011100110001100" OR uut_a_5_4 /= "111111101100011011100011110" OR uut_a_5_5 /= "000000011011100010101100100" THEN
              FAIL <= '1';
              FAIL_NUM <= "10000111";
              state <= "11111101";
            ELSE
              state <= "10010101";
            END IF;
            uut_rst <= '0';
          WHEN "10010101" =>
            uut_coord_shift <= "0110";
            uut_x <= "000000111000";
            uut_y <= "111110000101";
            uut_fx <= "0010110011";
            uut_fy <= "1111000001";
            uut_ft <= "1111000000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000001101010111100100000" OR uut_a_0_1 /= "000101110110010011110000000" OR uut_a_0_2 /= "000000101000000110101100000" OR uut_a_0_3 /= "000000000100100000110110000" OR uut_a_0_4 /= "000001111110010111101000000" OR uut_a_0_5 /= "000000001101100010100010000" OR uut_a_1_0 /= "000000001011101100100111100" OR uut_a_1_1 /= "000101000111100001010010000" OR uut_a_1_2 /= "000000100011000101110110100" OR uut_a_1_3 /= "000000000011111100101111010" OR uut_a_1_4 /= "000001101110100100101011000" OR uut_a_1_5 /= "000000001011110110001101110" OR uut_a_2_0 /= "000000000001010000001101011" OR uut_a_2_1 /= "000000100011000101110110100" OR uut_a_2_2 /= "000000000011110000101000001" OR uut_a_2_3 /= "000000000000011011000101000" OR uut_a_2_4 /= "000000001011110110001101110" OR uut_a_2_5 /= "000000000001010001001111001" OR uut_a_3_0 /= "000000000100100000110110000" OR uut_a_3_1 /= "000001111110010111101000000" OR uut_a_3_2 /= "000000001101100010100010000" OR uut_a_3_3 /= "000000000001100001100001000" OR uut_a_3_4 /= "000000101010101010011100000" OR uut_a_3_5 /= "000000000100100100100011000" OR uut_a_4_0 /= "000000000011111100101111010" OR uut_a_4_1 /= "000001101110100100101011000" OR uut_a_4_2 /= "000000001011110110001101110" OR uut_a_4_3 /= "000000000001010101010100111" OR uut_a_4_4 /= "000000100101010101001000100" OR uut_a_4_5 /= "000000000011111111111110101" OR uut_a_5_0 /= "000000000000011011000101000" OR uut_a_5_1 /= "000000001011110110001101110" OR uut_a_5_2 /= "000000000001010001001111001" OR uut_a_5_3 /= "000000000000001001001001000" OR uut_a_5_4 /= "000000000011111111111110101" OR uut_a_5_5 /= "000000000000011011011011010" THEN
              FAIL <= '1';
              FAIL_NUM <= "10001000";
              state <= "11111101";
            ELSE
              state <= "10010110";
            END IF;
            uut_rst <= '0';
          WHEN "10010110" =>
            uut_coord_shift <= "0110";
            uut_x <= "111110011110";
            uut_y <= "000001010000";
            uut_fx <= "1101001101";
            uut_fy <= "1011111100";
            uut_ft <= "1101011111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000111100100000" OR uut_a_0_1 /= "111111111111101001010100000" OR uut_a_0_2 /= "000000000001000100000100000" OR uut_a_0_3 /= "111111111111010010111110000" OR uut_a_0_4 /= "000000000010000111000110000" OR uut_a_0_5 /= "111111111001101010101110000" OR uut_a_1_0 /= "111111111111111111010010101" OR uut_a_1_1 /= "000000000000000010001000001" OR uut_a_1_2 /= "111111111111111001100111101" OR uut_a_1_3 /= "000000000000000100001110001" OR uut_a_1_4 /= "111111111111110011010101011" OR uut_a_1_5 /= "000000000000100101111111101" OR uut_a_2_0 /= "000000000000000010001000001" OR uut_a_2_1 /= "111111111111111001100111101" OR uut_a_2_2 /= "000000000000010011001001001" OR uut_a_2_3 /= "111111111111110011010101011" OR uut_a_2_4 /= "000000000000100101111111101" OR uut_a_2_5 /= "111111111110001110000000111" OR uut_a_3_0 /= "111111111111010010111110000" OR uut_a_3_1 /= "000000000010000111000110000" OR uut_a_3_2 /= "111111111001101010101110000" OR uut_a_3_3 /= "000000000100001100001001000" OR uut_a_3_4 /= "111111110011011011100101000" OR uut_a_3_5 /= "000000100101101101010001000" OR uut_a_4_0 /= "000000000000000100001110001" OR uut_a_4_1 /= "111111111111110011010101011" OR uut_a_4_2 /= "000000000000100101111111101" OR uut_a_4_3 /= "111111111111100110110111001" OR uut_a_4_4 /= "000000000001001011011010100" OR uut_a_4_5 /= "111111111100011101110000011" OR uut_a_5_0 /= "111111111111110011010101011" OR uut_a_5_1 /= "000000000000100101111111101" OR uut_a_5_2 /= "111111111110001110000000111" OR uut_a_5_3 /= "000000000001001011011010100" OR uut_a_5_4 /= "111111111100011101110000011" OR uut_a_5_5 /= "000000001010100110101110110" THEN
              FAIL <= '1';
              FAIL_NUM <= "10001001";
              state <= "11111101";
            ELSE
              state <= "10010111";
            END IF;
            uut_rst <= '0';
          WHEN "10010111" =>
            uut_coord_shift <= "0110";
            uut_x <= "111111100001";
            uut_y <= "000000001011";
            uut_fx <= "0000111111";
            uut_fy <= "1110010101";
            uut_ft <= "1110011000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000100001100001001000" OR uut_a_0_1 /= "000001010111111110111101000" OR uut_a_0_2 /= "000001011100001011000110000" OR uut_a_0_3 /= "111111111100111101100011000" OR uut_a_0_4 /= "111111000000001100011111000" OR uut_a_0_5 /= "111110111101001010000010000" OR uut_a_1_0 /= "000000000010101111111101111" OR uut_a_1_1 /= "000000111001101111010100000" OR uut_a_1_2 /= "000000111100011111010001111" OR uut_a_1_3 /= "111111111110000000011000111" OR uut_a_1_4 /= "111111010110001000001100010" OR uut_a_1_5 /= "111111010100001000100101010" OR uut_a_2_0 /= "000000000010111000010110001" OR uut_a_2_1 /= "000000111100011111010001111" OR uut_a_2_2 /= "000000111111010111101000001" OR uut_a_2_3 /= "111111111101111010010100000" OR uut_a_2_4 /= "111111010100001000100101010" OR uut_a_2_5 /= "111111010010000010111001011" OR uut_a_3_0 /= "111111111100111101100011000" OR uut_a_3_1 /= "111111000000001100011111000" OR uut_a_3_2 /= "111110111101001010000010000" OR uut_a_3_3 /= "000000000010001101000001000" OR uut_a_3_4 /= "000000101110010001010101000" OR uut_a_3_5 /= "000000110000011110010110000" OR uut_a_4_0 /= "111111111110000000011000111" OR uut_a_4_1 /= "111111010110001000001100010" OR uut_a_4_2 /= "111111010100001000100101010" OR uut_a_4_3 /= "000000000001011100100010101" OR uut_a_4_4 /= "000000011110010111010111110" OR uut_a_4_5 /= "000000011111110011111010011" OR uut_a_5_0 /= "111111111101111010010100000" OR uut_a_5_1 /= "111111010100001000100101010" OR uut_a_5_2 /= "111111010010000010111001011" OR uut_a_5_3 /= "000000000001100000111100101" OR uut_a_5_4 /= "000000011111110011111010011" OR uut_a_5_5 /= "000000100001010100110111001" THEN
              FAIL <= '1';
              FAIL_NUM <= "10001010";
              state <= "11111101";
            ELSE
              state <= "10011000";
            END IF;
            uut_rst <= '0';
          WHEN "10011000" =>
            uut_coord_shift <= "0110";
            uut_x <= "000000000011";
            uut_y <= "000000101000";
            uut_fx <= "0111001110";
            uut_fy <= "0011100100";
            uut_ft <= "1110011010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000010101111110010000000" OR uut_a_0_1 /= "001001011100001111111000000" OR uut_a_0_2 /= "000011100110101101101000000" OR uut_a_0_3 /= "111111110100011011011000000" OR uut_a_0_4 /= "111011000001110000110100000" OR uut_a_0_5 /= "111110000110011111011100000" OR uut_a_1_0 /= "000000010010111000011111110" OR uut_a_1_1 /= "001000000111010001101001001" OR uut_a_1_2 /= "000011000110010001001101011" OR uut_a_1_3 /= "111111110110000011100001101" OR uut_a_1_4 /= "111011101110100000111100101" OR uut_a_1_5 /= "111110010111100101000001000" OR uut_a_2_0 /= "000000000111001101011011010" OR uut_a_2_1 /= "000011000110010001001101011" OR uut_a_2_2 /= "000001001011101100111110001" OR uut_a_2_3 /= "111111111100001100111110111" OR uut_a_2_4 /= "111110010111100101000001000" OR uut_a_2_5 /= "111111011000001000010100001" OR uut_a_3_0 /= "111111110100011011011000000" OR uut_a_3_1 /= "111011000001110000110100000" OR uut_a_3_2 /= "111110000110011111011100000" OR uut_a_3_3 /= "000000000110000110000100000" OR uut_a_3_4 /= "000010100111100110101110000" OR uut_a_3_5 /= "000000111111111111101010000" OR uut_a_4_0 /= "111111110110000011100001101" OR uut_a_4_1 /= "111011101110100000111100101" OR uut_a_4_2 /= "111110010111100101000001000" OR uut_a_4_3 /= "000000000101001111001101011" OR uut_a_4_4 /= "000010010000000010010001100" OR uut_a_4_5 /= "000000110110111111101101000" OR uut_a_5_0 /= "111111111100001100111110111" OR uut_a_5_1 /= "111110010111100101000001000" OR uut_a_5_2 /= "111111011000001000010100001" OR uut_a_5_3 /= "000000000001111111111111010" OR uut_a_5_4 /= "000000110110111111101101000" OR uut_a_5_5 /= "000000010100111111111000110" THEN
              FAIL <= '1';
              FAIL_NUM <= "10001011";
              state <= "11111101";
            ELSE
              state <= "10011001";
            END IF;
            uut_rst <= '0';
          WHEN "10011001" =>
            uut_coord_shift <= "0110";
            uut_x <= "000001010100";
            uut_y <= "111110100011";
            uut_fx <= "1000111110";
            uut_fy <= "1001010110";
            uut_ft <= "1010101000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000011000000100001000000" OR uut_a_0_1 /= "111011101011010000100100000" OR uut_a_0_2 /= "000111111001010110101000000" OR uut_a_0_3 /= "000000010001001111000100000" OR uut_a_0_4 /= "111100111001110010110010000" OR uut_a_0_5 /= "000101101001111100010100000" OR uut_a_1_0 /= "111111111011101011010000100" OR uut_a_1_1 /= "000000110001101110100001100" OR uut_a_1_2 /= "111110100101001100011011110" OR uut_a_1_3 /= "111111111100111001110010110" OR uut_a_1_4 /= "000000100011100111011000000" OR uut_a_1_5 /= "111110111110111101101010011" OR uut_a_2_0 /= "000000000111111001010110101" OR uut_a_2_1 /= "111110100101001100011011110" OR uut_a_2_2 /= "000010100101110100011011001" OR uut_a_2_3 /= "000000000101101001111100010" OR uut_a_2_4 /= "111110111110111101101010011" OR uut_a_2_5 /= "000001110110110000110010100" OR uut_a_3_0 /= "000000010001001111000100000" OR uut_a_3_1 /= "111100111001110010110010000" OR uut_a_3_2 /= "000101101001111100010100000" OR uut_a_3_3 /= "000000001100010110000010000" OR uut_a_3_4 /= "111101110010000010101001000" OR uut_a_3_5 /= "000100000011001110101010000" OR uut_a_4_0 /= "111111111100111001110010110" OR uut_a_4_1 /= "000000100011100111011000000" OR uut_a_4_2 /= "111110111110111101101010011" OR uut_a_4_3 /= "111111111101110010000010101" OR uut_a_4_4 /= "000000011001100000100001101" OR uut_a_4_5 /= "111111010001011010110111011" OR uut_a_5_0 /= "000000000101101001111100010" OR uut_a_5_1 /= "111110111110111101101010011" OR uut_a_5_2 /= "000001110110110000110010100" OR uut_a_5_3 /= "000000000100000011001110101" OR uut_a_5_4 /= "111111010001011010110111011" OR uut_a_5_5 /= "000001010101000011110011110" THEN
              FAIL <= '1';
              FAIL_NUM <= "10001100";
              state <= "11111101";
            ELSE
              state <= "10011010";
            END IF;
            uut_rst <= '0';
          WHEN "10011010" =>
            uut_coord_shift <= "0110";
            uut_x <= "111111010100";
            uut_y <= "111111001110";
            uut_fx <= "1000001100";
            uut_fy <= "0000101001";
            uut_ft <= "1001100010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000011100011110100100100" OR uut_a_0_1 /= "001110011101100001100010010" OR uut_a_0_2 /= "111011010100111111000000110" OR uut_a_0_3 /= "000000011101011110101110000" OR uut_a_0_4 /= "001110111110000110010111000" OR uut_a_0_5 /= "111011001010011101011101000" OR uut_a_1_0 /= "000000001110011101100001100" OR uut_a_1_1 /= "000111010101111111100001111" OR uut_a_1_2 /= "111101101000001001111111111" OR uut_a_1_3 /= "000000001110111110000110010" OR uut_a_1_4 /= "000111100110100010001110101" OR uut_a_1_5 /= "111101100010110011111101001" OR uut_a_2_0 /= "111111111011010100111111000" OR uut_a_2_1 /= "111101101000001001111111111" OR uut_a_2_2 /= "000000110001000011101010011" OR uut_a_2_3 /= "111111111011001010011101011" OR uut_a_2_4 /= "111101100010110011111101001" OR uut_a_2_5 /= "000000110010110010001010101" OR uut_a_3_0 /= "000000011101011110101110000" OR uut_a_3_1 /= "001110111110000110010111000" OR uut_a_3_2 /= "111011001010011101011101000" OR uut_a_3_3 /= "000000011110100001001000000" OR uut_a_3_4 /= "001111011111110100100100000" OR uut_a_3_5 /= "111010111111100100001100000" OR uut_a_4_0 /= "000000001110111110000110010" OR uut_a_4_1 /= "000111100110100010001110101" OR uut_a_4_2 /= "111101100010110011111101001" OR uut_a_4_3 /= "000000001111011111110100100" OR uut_a_4_4 /= "000111110111101010001100010" OR uut_a_4_5 /= "111101011101010001111000000" OR uut_a_5_0 /= "111111111011001010011101011" OR uut_a_5_1 /= "111101100010110011111101001" OR uut_a_5_2 /= "000000110010110010001010101" OR uut_a_5_3 /= "111111111010111111100100001" OR uut_a_5_4 /= "111101011101010001111000000" OR uut_a_5_5 /= "000000110100100100100100000" THEN
              FAIL <= '1';
              FAIL_NUM <= "10001101";
              state <= "11111101";
            ELSE
              state <= "10011011";
            END IF;
            uut_rst <= '0';
          WHEN "10011011" =>
            uut_coord_shift <= "0110";
            uut_x <= "111110100110";
            uut_y <= "000000100001";
            uut_fx <= "0101110000";
            uut_fy <= "0111100110";
            uut_ft <= "0001001001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000001000001100000100100" OR uut_a_0_1 /= "111110001101010111000001000" OR uut_a_0_2 /= "111111010010111101100111010" OR uut_a_0_3 /= "111111110110110011001011100" OR uut_a_0_4 /= "000010000000110011011111000" OR uut_a_0_5 /= "000000110010100110100000110" OR uut_a_1_0 /= "111111111110001101010111000" OR uut_a_1_1 /= "000000011001000100111101110" OR uut_a_1_2 /= "000000001001110110100001011" OR uut_a_1_3 /= "000000000010000000110011011" OR uut_a_1_4 /= "111111100011110100101111001" OR uut_a_1_5 /= "111111110100111011100100110" OR uut_a_2_0 /= "111111111111010010111101100" OR uut_a_2_1 /= "000000001001110110100001011" OR uut_a_2_2 /= "000000000011110111101101001" OR uut_a_2_3 /= "000000000000110010100110100" OR uut_a_2_4 /= "111111110100111011100100110" OR uut_a_2_5 /= "111111111011101001101100001" OR uut_a_3_0 /= "111111110110110011001011100" OR uut_a_3_1 /= "000010000000110011011111000" OR uut_a_3_2 /= "000000110010100110100000110" OR uut_a_3_3 /= "000000001010010101100100100" OR uut_a_3_4 /= "111101101111010010000001000" OR uut_a_3_5 /= "111111000111001001010111010" OR uut_a_4_0 /= "000000000010000000110011011" OR uut_a_4_1 /= "111111100011110100101111001" OR uut_a_4_2 /= "111111110100111011100100110" OR uut_a_4_3 /= "111111111101101111010010000" OR uut_a_4_4 /= "000000011111101010000011110" OR uut_a_4_5 /= "000000001100011011111100111" OR uut_a_5_0 /= "000000000000110010100110100" OR uut_a_5_1 /= "111111110100111011100100110" OR uut_a_5_2 /= "111111111011101001101100001" OR uut_a_5_3 /= "111111111111000111001001010" OR uut_a_5_4 /= "000000001100011011111100111" OR uut_a_5_5 /= "000000000100111000101100100" THEN
              FAIL <= '1';
              FAIL_NUM <= "10001110";
              state <= "11111101";
            ELSE
              state <= "10011100";
            END IF;
            uut_rst <= '0';
          WHEN "10011100" =>
            uut_coord_shift <= "0110";
            uut_x <= "000001111111";
            uut_y <= "000000001101";
            uut_fx <= "0000010000";
            uut_fy <= "1101010011";
            uut_ft <= "1110111000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001001111101100100" OR uut_a_0_1 /= "000001000001011000000000010" OR uut_a_0_2 /= "000000001000101101110111100" OR uut_a_0_3 /= "111111111011100011111100000" OR uut_a_0_4 /= "111100010110111110101110000" OR uut_a_0_5 /= "111111100000111011100100000" OR uut_a_1_0 /= "000000000001000001011000000" OR uut_a_1_1 /= "000000110101101000001100001" OR uut_a_1_2 /= "000000000111001001101000000" OR uut_a_1_3 /= "111111111100010110111110101" OR uut_a_1_4 /= "111101000000110110011100101" OR uut_a_1_5 /= "111111100110100000110111000" OR uut_a_2_0 /= "000000000000001000101101110" OR uut_a_2_1 /= "000000000111001001101000000" OR uut_a_2_2 /= "000000000000111101000001000" OR uut_a_2_3 /= "111111111111100000111011100" OR uut_a_2_4 /= "111111100110100000110111000" OR uut_a_2_5 /= "111111111100100110100000111" OR uut_a_3_0 /= "111111111011100011111100000" OR uut_a_3_1 /= "111100010110111110101110000" OR uut_a_3_2 /= "111111100000111011100100000" OR uut_a_3_3 /= "000000001111110100100000000" OR uut_a_3_4 /= "001100111110100100010000000" OR uut_a_3_5 /= "000001101110101111100000000" OR uut_a_4_0 /= "111111111100010110111110101" OR uut_a_4_1 /= "111101000000110110011100101" OR uut_a_4_2 /= "111111100110100000110111000" OR uut_a_4_3 /= "000000001100111110100100010" OR uut_a_4_4 /= "001010101001010100101111001" OR uut_a_4_5 /= "000001011010110101111101110" OR uut_a_5_0 /= "111111111111100000111011100" OR uut_a_5_1 /= "111111100110100000110111000" OR uut_a_5_2 /= "111111111100100110100000111" OR uut_a_5_3 /= "000000000001101110101111100" OR uut_a_5_4 /= "000001011010110101111101110" OR uut_a_5_5 /= "000000001100000111001100100" THEN
              FAIL <= '1';
              FAIL_NUM <= "10001111";
              state <= "11111101";
            ELSE
              state <= "10011101";
            END IF;
            uut_rst <= '0';
          WHEN "10011101" =>
            uut_coord_shift <= "0110";
            uut_x <= "111111111110";
            uut_y <= "111110010011";
            uut_fx <= "0110001101";
            uut_fy <= "1001000010";
            uut_ft <= "1110111111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000010100011010111000100" OR uut_a_0_1 /= "111110000101011110101101000" OR uut_a_0_2 /= "110100000010001111111001010" OR uut_a_0_3 /= "000000001101011011100010100" OR uut_a_0_4 /= "111110101111011010110001000" OR uut_a_0_5 /= "111000001000010111010010010" OR uut_a_1_0 /= "111111111110000101011110101" OR uut_a_1_1 /= "000000001011011111000111110" OR uut_a_1_2 /= "000001000111110010100000101" OR uut_a_1_3 /= "111111111110101111011010110" OR uut_a_1_4 /= "000000000111100011011111011" OR uut_a_1_5 /= "000000101111001101110100010" OR uut_a_2_0 /= "111111110100000010001111111" OR uut_a_2_1 /= "000001000111110010100000101" OR uut_a_2_2 /= "000111000000101011101011111" OR uut_a_2_3 /= "111111111000001000010111010" OR uut_a_2_4 /= "000000101111001101110100010" OR uut_a_2_5 /= "000100100111000110010110110" OR uut_a_3_0 /= "000000001101011011100010100" OR uut_a_3_1 /= "111110101111011010110001000" OR uut_a_3_2 /= "111000001000010111010010010" OR uut_a_3_3 /= "000000001000110101010100100" OR uut_a_3_4 /= "111111001011000000000101000" OR uut_a_3_5 /= "111010110100110000011111010" OR uut_a_4_0 /= "111111111110101111011010110" OR uut_a_4_1 /= "000000000111100011011111011" OR uut_a_4_2 /= "000000101111001101110100010" OR uut_a_4_3 /= "111111111111001011000000000" OR uut_a_4_4 /= "000000000100111101111111100" OR uut_a_4_5 /= "000000011111000011011101000" OR uut_a_5_0 /= "111111111000001000010111010" OR uut_a_5_1 /= "000000101111001101110100010" OR uut_a_5_2 /= "000100100111000110010110110" OR uut_a_5_3 /= "111111111010110100110000011" OR uut_a_5_4 /= "000000011111000011011101000" OR uut_a_5_5 /= "000011000010000101100101101" THEN
              FAIL <= '1';
              FAIL_NUM <= "10010000";
              state <= "11111101";
            ELSE
              state <= "10011110";
            END IF;
            uut_rst <= '0';
          WHEN "10011110" =>
            uut_coord_shift <= "0110";
            uut_x <= "000001010011";
            uut_y <= "111111100110";
            uut_fx <= "0001110100";
            uut_fy <= "0101000110";
            uut_ft <= "0110001100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000011011100100000000" OR uut_a_0_1 /= "111110100001010000010000000" OR uut_a_0_2 /= "000001001011110011000000000" OR uut_a_0_3 /= "111111111000000101011000000" OR uut_a_0_4 /= "000011011001101100001100000" OR uut_a_0_5 /= "111101010001110110010000000" OR uut_a_1_0 /= "111111111110100001010000010" OR uut_a_1_1 /= "000000101000101101100001001" OR uut_a_1_2 /= "111111011111011011100101100" OR uut_a_1_3 /= "000000000011011001101100001" OR uut_a_1_4 /= "111110100010011101100000110" OR uut_a_1_5 /= "000001001010110101001100001" OR uut_a_2_0 /= "000000000001001011110011000" OR uut_a_2_1 /= "111111011111011011100101100" OR uut_a_2_2 /= "000000011010000011100010000" OR uut_a_2_3 /= "111111111101010001110110010" OR uut_a_2_4 /= "000001001010110101001100001" OR uut_a_2_5 /= "111111000100001000101001100" OR uut_a_3_0 /= "111111111000000101011000000" OR uut_a_3_1 /= "000011011001101100001100000" OR uut_a_3_2 /= "111101010001110110010000000" OR uut_a_3_3 /= "000000010010001100000010000" OR uut_a_3_4 /= "111000001011110101001001000" OR uut_a_3_5 /= "000110010000001000101100000" OR uut_a_4_0 /= "000000000011011001101100001" OR uut_a_4_1 /= "111110100010011101100000110" OR uut_a_4_2 /= "000001001010110101001100001" OR uut_a_4_3 /= "111111111000001011110101001" OR uut_a_4_4 /= "000011010110111010101010101" OR uut_a_4_5 /= "111101010100000100010001000" OR uut_a_5_0 /= "111111111101010001110110010" OR uut_a_5_1 /= "000001001010110101001100001" OR uut_a_5_2 /= "111111000100001000101001100" OR uut_a_5_3 /= "000000000110010000001000101" OR uut_a_5_4 /= "111101010100000100010001000" OR uut_a_5_5 /= "000010001001100010111111001" THEN
              FAIL <= '1';
              FAIL_NUM <= "10010001";
              state <= "11111101";
            ELSE
              state <= "10011111";
            END IF;
            uut_rst <= '0';
          WHEN "10011111" =>
            uut_coord_shift <= "0110";
            uut_x <= "000001101110";
            uut_y <= "111110110001";
            uut_fx <= "1100001001";
            uut_fy <= "0110010111";
            uut_ft <= "0001100000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000110000001000010000" OR uut_a_0_1 /= "111101010100100010100111000" OR uut_a_0_2 /= "000010100101011100010111000" OR uut_a_0_3 /= "111111110100111111110110000" OR uut_a_0_4 /= "000100111001100100011101000" OR uut_a_0_5 /= "111011010001011011101101000" OR uut_a_1_0 /= "111111111101010100100010100" OR uut_a_1_1 /= "000001001100010110100101101" OR uut_a_1_2 /= "111110110110010100110111110" OR uut_a_1_3 /= "000000000100111001100100011" OR uut_a_1_4 /= "111101110100010111010001000" OR uut_a_1_5 /= "000010000110101111001010011" OR uut_a_2_0 /= "000000000010100101011100010" OR uut_a_2_1 /= "111110110110010100110111110" OR uut_a_2_2 /= "000001000111000101101011111" OR uut_a_2_3 /= "111111111011010001011011101" OR uut_a_2_4 /= "000010000110101111001010011" OR uut_a_2_5 /= "111101111101111111011001110" OR uut_a_3_0 /= "111111110100111111110110000" OR uut_a_3_1 /= "000100111001100100011101000" OR uut_a_3_2 /= "111011010001011011101101000" OR uut_a_3_3 /= "000000010100000111110010000" OR uut_a_3_4 /= "110111000010100010001111000" OR uut_a_3_5 /= "001000101001010101111111000" OR uut_a_4_0 /= "000000000100111001100100011" OR uut_a_4_1 /= "111101110100010111010001000" OR uut_a_4_2 /= "000010000110101111001010011" OR uut_a_4_3 /= "111111110111000010100010001" OR uut_a_4_4 /= "000011111111010111110000010" OR uut_a_4_5 /= "111100001001100101101101011" OR uut_a_5_0 /= "111111111011010001011011101" OR uut_a_5_1 /= "000010000110101111001010011" OR uut_a_5_2 /= "111101111101111111011001110" OR uut_a_5_3 /= "000000001000101001010101111" OR uut_a_5_4 /= "111100001001100101101101011" OR uut_a_5_5 /= "000011101101110000111100100" THEN
              FAIL <= '1';
              FAIL_NUM <= "10010010";
              state <= "11111101";
            ELSE
              state <= "10100000";
            END IF;
            uut_rst <= '0';
          WHEN "10100000" =>
            uut_coord_shift <= "0111";
            uut_x <= "000000000001";
            uut_y <= "000000111001";
            uut_fx <= "0101000111";
            uut_fy <= "0000100001";
            uut_ft <= "1011001111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000100110101011000100" OR uut_a_0_1 /= "111110111100010100101001000" OR uut_a_0_2 /= "000000000000000000000000000" OR uut_a_0_3 /= "000000001000010011101101000" OR uut_a_0_4 /= "111110001011101100001010000" OR uut_a_0_5 /= "000000000000000000000000000" OR uut_a_1_0 /= "111111111110111100010100101" OR uut_a_1_1 /= "000000001110110011011111000" OR uut_a_1_2 /= "000000000000000000000000000" OR uut_a_1_3 /= "111111111110001011101100001" OR uut_a_1_4 /= "000000011001011100010101110" OR uut_a_1_5 /= "000000000000000000000000000" OR uut_a_2_0 /= "000000000000000000000000000" OR uut_a_2_1 /= "000000000000000000000000000" OR uut_a_2_2 /= "000000000000000000000000000" OR uut_a_2_3 /= "000000000000000000000000000" OR uut_a_2_4 /= "000000000000000000000000000" OR uut_a_2_5 /= "000000000000000000000000000" OR uut_a_3_0 /= "000000001000010011101101000" OR uut_a_3_1 /= "111110001011101100001010000" OR uut_a_3_2 /= "000000000000000000000000000" OR uut_a_3_3 /= "000000001110010001110010000" OR uut_a_3_4 /= "111100111000000111000100000" OR uut_a_3_5 /= "000000000000000000000000000" OR uut_a_4_0 /= "111111111110001011101100001" OR uut_a_4_1 /= "000000011001011100010101110" OR uut_a_4_2 /= "000000000000000000000000000" OR uut_a_4_3 /= "111111111100111000000111000" OR uut_a_4_4 /= "000000101011101110011101001" OR uut_a_4_5 /= "000000000000000000000000000" OR uut_a_5_0 /= "000000000000000000000000000" OR uut_a_5_1 /= "000000000000000000000000000" OR uut_a_5_2 /= "000000000000000000000000000" OR uut_a_5_3 /= "000000000000000000000000000" OR uut_a_5_4 /= "000000000000000000000000000" OR uut_a_5_5 /= "000000000000000000000000000" THEN
              FAIL <= '1';
              FAIL_NUM <= "10010011";
              state <= "11111101";
            ELSE
              state <= "10100001";
            END IF;
            uut_rst <= '0';
          WHEN "10100001" =>
            uut_coord_shift <= "0111";
            uut_x <= "111111101001";
            uut_y <= "111111011100";
            uut_fx <= "0111011101";
            uut_fy <= "0001111011";
            uut_ft <= "0011001000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000001111110100100" OR uut_a_0_1 /= "000000000010010110010010110" OR uut_a_0_2 /= "111111111010100011111101000" OR uut_a_0_3 /= "111111111110110011000000100" OR uut_a_0_4 /= "111111110100100100100100110" OR uut_a_0_5 /= "000000011010011101110101000" OR uut_a_1_0 /= "000000000000000010010110010" OR uut_a_1_1 /= "000000000000010110010011110" OR uut_a_1_2 /= "111111111111001100010101100" OR uut_a_1_3 /= "111111111111110100100100100" OR uut_a_1_4 /= "111111111110010011011011011" OR uut_a_1_5 /= "000000000011111011011011010" OR uut_a_2_0 /= "111111111111111010100011111" OR uut_a_2_1 /= "111111111111001100010101100" OR uut_a_2_2 /= "000000000001110111101001000" OR uut_a_2_3 /= "000000000000011010011101110" OR uut_a_2_4 /= "000000000011111011011011010" OR uut_a_2_5 /= "111111110110111001101111110" OR uut_a_3_0 /= "111111111110110011000000100" OR uut_a_3_1 /= "111111110100100100100100110" OR uut_a_3_2 /= "000000011010011101110101000" OR uut_a_3_3 /= "000000000101110110101100100" OR uut_a_3_4 /= "000000110111100111100110110" OR uut_a_3_5 /= "111101111111001100101101000" OR uut_a_4_0 /= "111111111111110100100100100" OR uut_a_4_1 /= "111111111110010011011011011" OR uut_a_4_2 /= "000000000011111011011011010" OR uut_a_4_3 /= "000000000000110111100111100" OR uut_a_4_4 /= "000000001000010000011000010" OR uut_a_4_5 /= "111111101100111000011000101" OR uut_a_5_0 /= "000000000000011010011101110" OR uut_a_5_1 /= "000000000011111011011011010" OR uut_a_5_2 /= "111111110110111001101111110" OR uut_a_5_3 /= "111111111101111111001100101" OR uut_a_5_4 /= "111111101100111000011000101" OR uut_a_5_5 /= "000000101100010001101000100" THEN
              FAIL <= '1';
              FAIL_NUM <= "10010100";
              state <= "11111101";
            ELSE
              state <= "10100010";
            END IF;
            uut_rst <= '0';
          WHEN "10100010" =>
            uut_coord_shift <= "0111";
            uut_x <= "000001110000";
            uut_y <= "111110110010";
            uut_fx <= "0000010001";
            uut_fy <= "0000111010";
            uut_ft <= "1010100000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000011111010010100100" OR uut_a_0_1 /= "000001101101100000111110000" OR uut_a_0_2 /= "111100001111011101010011010" OR uut_a_0_3 /= "111111111110100111111001100" OR uut_a_0_4 /= "111111011001011101001010000" OR uut_a_0_5 /= "000001010100101010001111110" OR uut_a_1_0 /= "000000000001101101100000111" OR uut_a_1_1 /= "000000101111111010011011001" OR uut_a_1_2 /= "111110010110110000110100011" OR uut_a_1_3 /= "111111111111011001011101001" OR uut_a_1_4 /= "111111101111001000110000011" OR uut_a_1_5 /= "000000100101000010011110111" OR uut_a_2_0 /= "111111111100001111011101010" OR uut_a_2_1 /= "111110010110110000110100011" OR uut_a_2_2 /= "000011100111001001010110000" OR uut_a_2_3 /= "000000000001010100101010001" OR uut_a_2_4 /= "000000100101000010011110111" OR uut_a_2_5 /= "111110101110101001011001110" OR uut_a_3_0 /= "111111111110100111111001100" OR uut_a_3_1 /= "111111011001011101001010000" OR uut_a_3_2 /= "000001010100101010001111110" OR uut_a_3_3 /= "000000000000011111000000100" OR uut_a_3_4 /= "000000001101100100001110000" OR uut_a_3_5 /= "111111100010001101000001010" OR uut_a_4_0 /= "111111111111011001011101001" OR uut_a_4_1 /= "111111101111001000110000011" OR uut_a_4_2 /= "000000100101000010011110111" OR uut_a_4_3 /= "000000000000001101100100001" OR uut_a_4_4 /= "000000000101111011110110001" OR uut_a_4_5 /= "111111110010111101101100100" OR uut_a_5_0 /= "000000000001010100101010001" OR uut_a_5_1 /= "000000100101000010011110111" OR uut_a_5_2 /= "111110101110101001011001110" OR uut_a_5_3 /= "111111111111100010001101000" OR uut_a_5_4 /= "111111110010111101101100100" OR uut_a_5_5 /= "000000011100101000011111010" THEN
              FAIL <= '1';
              FAIL_NUM <= "10010101";
              state <= "11111101";
            ELSE
              state <= "10100011";
            END IF;
            uut_rst <= '0';
          WHEN "10100011" =>
            uut_coord_shift <= "0111";
            uut_x <= "000000011111";
            uut_y <= "000001100011";
            uut_fx <= "1110110101";
            uut_fy <= "0101011000";
            uut_ft <= "0011101101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000011111010010100100" OR uut_a_0_1 /= "111101000000010110010011100" OR uut_a_0_2 /= "000010011100011100110100000" OR uut_a_0_3 /= "000000000101101011100110000" OR uut_a_0_4 /= "111011101001100111111010000" OR uut_a_0_5 /= "000011100011001111110000000" OR uut_a_1_0 /= "111111111101000000010110010" OR uut_a_1_1 /= "000010010010101110111011000" OR uut_a_1_2 /= "111110001000001101111100001" OR uut_a_1_3 /= "111111111011101001100111111" OR uut_a_1_4 /= "000011010101001000011100100" OR uut_a_1_5 /= "111101010010000000111100010" OR uut_a_2_0 /= "000000000010011100011100110" OR uut_a_2_1 /= "111110001000001101111100001" OR uut_a_2_2 /= "000001100001110010000000100" OR uut_a_2_3 /= "000000000011100011001111110" OR uut_a_2_4 /= "111101010010000000111100010" OR uut_a_2_5 /= "000010001110000001110110000" OR uut_a_3_0 /= "000000000101101011100110000" OR uut_a_3_1 /= "111011101001100111111010000" OR uut_a_3_2 /= "000011100011001111110000000" OR uut_a_3_3 /= "000000001000010000001000000" OR uut_a_3_4 /= "111001101011101001111000000" OR uut_a_3_5 /= "000101001010000101000000000" OR uut_a_4_0 /= "111111111011101001100111111" OR uut_a_4_1 /= "000011010101001000011100100" OR uut_a_4_2 /= "111101010010000000111100010" OR uut_a_4_3 /= "111111111001101011101001111" OR uut_a_4_4 /= "000100110101100100111100001" OR uut_a_4_5 /= "111100000011010010001011000" OR uut_a_5_0 /= "000000000011100011001111110" OR uut_a_5_1 /= "111101010010000000111100010" OR uut_a_5_2 /= "000010001110000001110110000" OR uut_a_5_3 /= "000000000101001010000101000" OR uut_a_5_4 /= "111100000011010010001011000" OR uut_a_5_5 /= "000011001110010011001000000" THEN
              FAIL <= '1';
              FAIL_NUM <= "10010110";
              state <= "11111101";
            ELSE
              state <= "10100100";
            END IF;
            uut_rst <= '0';
          WHEN "10100100" =>
            uut_coord_shift <= "0111";
            uut_x <= "111110111001";
            uut_y <= "111111101001";
            uut_fx <= "1110001100";
            uut_fy <= "0100011010";
            uut_ft <= "0011110000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000011111000000100" OR uut_a_0_1 /= "111111111000011111011000010" OR uut_a_0_2 /= "000000000010101010100010110" OR uut_a_0_3 /= "111111111111001011010101100" OR uut_a_0_4 /= "000000001100110000010010110" OR uut_a_0_5 /= "111111111011011110010110010" OR uut_a_1_0 /= "111111111111111000011111011" OR uut_a_1_1 /= "000000000001110100011001101" OR uut_a_1_2 /= "111111111111010110101100100" OR uut_a_1_3 /= "000000000000001100110000010" OR uut_a_1_4 /= "111111111100111010010011011" OR uut_a_1_5 /= "000000000001000110001001100" OR uut_a_2_0 /= "000000000000000010101010100" OR uut_a_2_1 /= "111111111111010110101100100" OR uut_a_2_2 /= "000000000000001110101001111" OR uut_a_2_3 /= "111111111111111011011110010" OR uut_a_2_4 /= "000000000001000110001001100" OR uut_a_2_5 /= "111111111111100111000110111" OR uut_a_3_0 /= "111111111111001011010101100" OR uut_a_3_1 /= "000000001100110000010010110" OR uut_a_3_2 /= "111111111011011110010110010" OR uut_a_3_3 /= "000000000001011001011100100" OR uut_a_3_4 /= "111111101010010101100110010" OR uut_a_3_5 /= "000000000111101011111100110" OR uut_a_4_0 /= "000000000000001100110000010" OR uut_a_4_1 /= "111111111100111010010011011" OR uut_a_4_2 /= "000000000001000110001001100" OR uut_a_4_3 /= "111111111111101010010101100" OR uut_a_4_4 /= "000000000101001111110001001" OR uut_a_4_5 /= "111111111110001000110110110" OR uut_a_5_0 /= "111111111111111011011110010" OR uut_a_5_1 /= "000000000001000110001001100" OR uut_a_5_2 /= "111111111111100111000110111" OR uut_a_5_3 /= "000000000000000111101011111" OR uut_a_5_4 /= "111111111110001000110110110" OR uut_a_5_5 /= "000000000000101010010001101" THEN
              FAIL <= '1';
              FAIL_NUM <= "10010111";
              state <= "11111101";
            ELSE
              state <= "10100101";
            END IF;
            uut_rst <= '0';
          WHEN "10100101" =>
            uut_coord_shift <= "0111";
            uut_x <= "111111011101";
            uut_y <= "000001100011";
            uut_fx <= "0111001000";
            uut_fy <= "0100100011";
            uut_ft <= "0011010011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000011010000011100010000" OR uut_a_0_1 /= "000000100111000101010011000" OR uut_a_0_2 /= "001000001001000110101000000" OR uut_a_0_3 /= "000000001100110110111100000" OR uut_a_0_4 /= "000000010011010010011010000" OR uut_a_0_5 /= "000100000001001010110000000" OR uut_a_1_0 /= "000000000000100111000101010" OR uut_a_1_1 /= "000000000000111010100111111" OR uut_a_1_2 /= "000000001100001101101001111" OR uut_a_1_3 /= "000000000000010011010010011" OR uut_a_1_4 /= "000000000000011100111011100" OR uut_a_1_5 /= "000000000110000001110000001" OR uut_a_2_0 /= "000000001000001001000110101" OR uut_a_2_1 /= "000000001100001101101001111" OR uut_a_2_2 /= "000010100010110110000100100" OR uut_a_2_3 /= "000000000100000001001010110" OR uut_a_2_4 /= "000000000110000001110000001" OR uut_a_2_5 /= "000001010000010111010111000" OR uut_a_3_0 /= "000000001100110110111100000" OR uut_a_3_1 /= "000000010011010010011010000" OR uut_a_3_2 /= "000100000001001010110000000" OR uut_a_3_3 /= "000000000110010110001000000" OR uut_a_3_4 /= "000000001001100001001100000" OR uut_a_3_5 /= "000001111110111010100000000" OR uut_a_4_0 /= "000000000000010011010010011" OR uut_a_4_1 /= "000000000000011100111011100" OR uut_a_4_2 /= "000000000110000001110000001" OR uut_a_4_3 /= "000000000000001001100001001" OR uut_a_4_4 /= "000000000000001110010001110" OR uut_a_4_5 /= "000000000010111110010111110" OR uut_a_5_0 /= "000000000100000001001010110" OR uut_a_5_1 /= "000000000110000001110000001" OR uut_a_5_2 /= "000001010000010111010111000" OR uut_a_5_3 /= "000000000001111110111010100" OR uut_a_5_4 /= "000000000010111110010111110" OR uut_a_5_5 /= "000000100111101010010010000" THEN
              FAIL <= '1';
              FAIL_NUM <= "10011000";
              state <= "11111101";
            ELSE
              state <= "10100110";
            END IF;
            uut_rst <= '0';
          WHEN "10100110" =>
            uut_coord_shift <= "0111";
            uut_x <= "111100111000";
            uut_y <= "111111001000";
            uut_fx <= "0001011101";
            uut_fy <= "1111010110";
            uut_ft <= "1000110100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000011000101110000010000" OR uut_a_0_1 /= "010000001110001101010100000" OR uut_a_0_2 /= "101110000010100011100011000" OR uut_a_0_3 /= "000000010111011001101010000" OR uut_a_0_4 /= "001111010110110101100100000" OR uut_a_0_5 /= "101110111111110110111111000" OR uut_a_1_0 /= "000000010000001110001101010" OR uut_a_1_1 /= "001010101001010100101111001" OR uut_a_1_2 /= "110100001101101011010100111" OR uut_a_1_3 /= "000000001111010110110101100" OR uut_a_1_4 /= "001010000100111111001001101" OR uut_a_1_5 /= "110100110101111010000101010" OR uut_a_2_0 /= "111111101110000010100011100" OR uut_a_2_1 /= "110100001101101011010100111" OR uut_a_2_2 /= "001101000011001001001011000" OR uut_a_2_3 /= "111111101110111111110110111" OR uut_a_2_4 /= "110100110101111010000101010" OR uut_a_2_5 /= "001100010110100110100011001" OR uut_a_3_0 /= "000000010111011001101010000" OR uut_a_3_1 /= "001111010110110101100100000" OR uut_a_3_2 /= "101110111111110110111111000" OR uut_a_3_3 /= "000000010110001001110010000" OR uut_a_3_4 /= "001110100010011010110100000" OR uut_a_3_5 /= "101111111001111001001011000" OR uut_a_4_0 /= "000000001111010110110101100" OR uut_a_4_1 /= "001010000100111111001001101" OR uut_a_4_2 /= "110100110101111010000101010" OR uut_a_4_3 /= "000000001110100010011010110" OR uut_a_4_4 /= "001001100010100101100110001" OR uut_a_4_5 /= "110101011011111111100001001" OR uut_a_5_0 /= "111111101110111111110110111" OR uut_a_5_1 /= "110100110101111010000101010" OR uut_a_5_2 /= "001100010110100110100011001" OR uut_a_5_3 /= "111111101111111001111001001" OR uut_a_5_4 /= "110101011011111111100001001" OR uut_a_5_5 /= "001011101100011011111101100" THEN
              FAIL <= '1';
              FAIL_NUM <= "10011001";
              state <= "11111101";
            ELSE
              state <= "10100111";
            END IF;
            uut_rst <= '0';
          WHEN "10100111" =>
            uut_coord_shift <= "0111";
            uut_x <= "111101110110";
            uut_y <= "000010101011";
            uut_fx <= "1000010000";
            uut_fy <= "0101110100";
            uut_ft <= "1001010000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000011110100001001000000" OR uut_a_0_1 /= "110101100000100111010000000" OR uut_a_0_2 /= "110100000101000011111000000" OR uut_a_0_3 /= "111111111101011111110110000" OR uut_a_0_4 /= "000000110111000011011100000" OR uut_a_0_5 /= "000000111110100011111010000" OR uut_a_1_0 /= "111111110101100000100111010" OR uut_a_1_1 /= "000011100110110010100000100" OR uut_a_1_2 /= "000100000110010000101010110" OR uut_a_1_3 /= "000000000000110111000011011" OR uut_a_1_4 /= "111111101101000100110100011" OR uut_a_1_5 /= "111111101010011111101010000" OR uut_a_2_0 /= "111111110100000101000011111" OR uut_a_2_1 /= "000100000110010000101010110" OR uut_a_2_2 /= "000100101010000001011111001" OR uut_a_2_3 /= "000000000000111110100011111" OR uut_a_2_4 /= "111111101010011111101010000" OR uut_a_2_5 /= "111111100111100011111110010" OR uut_a_3_0 /= "111111111101011111110110000" OR uut_a_3_1 /= "000000110111000011011100000" OR uut_a_3_2 /= "000000111110100011111010000" OR uut_a_3_3 /= "000000000000001101001000100" OR uut_a_3_4 /= "111111111011011111000101000" OR uut_a_3_5 /= "111111111010110111101011100" OR uut_a_4_0 /= "000000000000110111000011011" OR uut_a_4_1 /= "111111101101000100110100011" OR uut_a_4_2 /= "111111101010011111101010000" OR uut_a_4_3 /= "111111111111111011011111000" OR uut_a_4_4 /= "000000000001100011010100010" OR uut_a_4_5 /= "000000000001110000110111000" OR uut_a_5_0 /= "000000000000111110100011111" OR uut_a_5_1 /= "111111101010011111101010000" OR uut_a_5_2 /= "111111100111100011111110010" OR uut_a_5_3 /= "111111111111111010110111101" OR uut_a_5_4 /= "000000000001110000110111000" OR uut_a_5_5 /= "000000000010000000010000000" THEN
              FAIL <= '1';
              FAIL_NUM <= "10011010";
              state <= "11111101";
            ELSE
              state <= "10101000";
            END IF;
            uut_rst <= '0';
          WHEN "10101000" =>
            uut_coord_shift <= "0111";
            uut_x <= "000001010110";
            uut_y <= "000000000000";
            uut_fx <= "1011011111";
            uut_fy <= "0001001001";
            uut_ft <= "1001111101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000010000100010000000000" OR uut_a_0_1 /= "110100011000000110000000000" OR uut_a_0_2 /= "000100010000110001000000000" OR uut_a_0_3 /= "000000010101110101010000000" OR uut_a_0_4 /= "110000101001100011110000000" OR uut_a_0_5 /= "000101101000001110101000000" OR uut_a_1_0 /= "111111110100011000000110000" OR uut_a_1_1 /= "001000001011000011110010000" OR uut_a_1_2 /= "111101000000001101100011000" OR uut_a_1_3 /= "111111110000101001100011110" OR uut_a_1_4 /= "001010110010110001110111010" OR uut_a_1_5 /= "111100000010101101101101111" OR uut_a_2_0 /= "000000000100010000110001000" OR uut_a_2_1 /= "111101000000001101100011000" OR uut_a_2_2 /= "000001000110010100101000100" OR uut_a_2_3 /= "000000000101101000001110101" OR uut_a_2_4 /= "111100000010101101101101111" OR uut_a_2_5 /= "000001011100110111110001010" OR uut_a_3_0 /= "000000010101110101010000000" OR uut_a_3_1 /= "110000101001100011110000000" OR uut_a_3_2 /= "000101101000001110101000000" OR uut_a_3_3 /= "000000011100110101010010000" OR uut_a_3_4 /= "101011101110100010010110000" OR uut_a_3_5 /= "000111011011101111001001000" OR uut_a_4_0 /= "111111110000101001100011110" OR uut_a_4_1 /= "001010110010110001110111010" OR uut_a_4_2 /= "111100000010101101101101111" OR uut_a_4_3 /= "111111101011101110100010010" OR uut_a_4_4 /= "001110010000010001110110100" OR uut_a_4_5 /= "111010110001011111110110101" OR uut_a_5_0 /= "000000000101101000001110101" OR uut_a_5_1 /= "111100000010101101101101111" OR uut_a_5_2 /= "000001011100110111110001010" OR uut_a_5_3 /= "000000000111011011101111001" OR uut_a_5_4 /= "111010110001011111110110101" OR uut_a_5_5 /= "000001111010101001101001110" THEN
              FAIL <= '1';
              FAIL_NUM <= "10011011";
              state <= "11111101";
            ELSE
              state <= "10101001";
            END IF;
            uut_rst <= '0';
          WHEN "10101001" =>
            uut_coord_shift <= "0111";
            uut_x <= "000001010111";
            uut_y <= "000000110010";
            uut_fx <= "1000111001";
            uut_fy <= "1000111010";
            uut_ft <= "1010011100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000010000000000" OR uut_a_0_1 /= "000000000001111111000000000" OR uut_a_0_2 /= "000000000000001101000000000" OR uut_a_0_3 /= "111111111111101010011000000" OR uut_a_0_4 /= "111111101010100010110100000" OR uut_a_0_5 /= "111111111101110011011100000" OR uut_a_1_0 /= "000000000000000001111111000" OR uut_a_1_1 /= "000000000001111110000000100" OR uut_a_1_2 /= "000000000000001100111001100" OR uut_a_1_3 /= "111111111111101010100010110" OR uut_a_1_4 /= "111111101010101101100010100" OR uut_a_1_5 /= "111111111101110100100010010" OR uut_a_2_0 /= "000000000000000000001101000" OR uut_a_2_1 /= "000000000000001100111001100" OR uut_a_2_2 /= "000000000000000001010100100" OR uut_a_2_3 /= "111111111111111101110011011" OR uut_a_2_4 /= "111111111101110100100010010" OR uut_a_2_5 /= "111111111111110001101110010" OR uut_a_3_0 /= "111111111111101010011000000" OR uut_a_3_1 /= "111111101010100010110100000" OR uut_a_3_2 /= "111111111101110011011100000" OR uut_a_3_3 /= "000000000011101001110100100" OR uut_a_3_4 /= "000011100111111111100101110" OR uut_a_3_5 /= "000000010111101111110101010" OR uut_a_4_0 /= "111111111111101010100010110" OR uut_a_4_1 /= "111111101010101101100010100" OR uut_a_4_2 /= "111111111101110100100010010" OR uut_a_4_3 /= "000000000011100111111111100" OR uut_a_4_4 /= "000011100110001011100101111" OR uut_a_4_5 /= "000000010111100011111101010" OR uut_a_5_0 /= "111111111111111101110011011" OR uut_a_5_1 /= "111111111101110100100010010" OR uut_a_5_2 /= "111111111111110001101110010" OR uut_a_5_3 /= "000000000000010111101111110" OR uut_a_5_4 /= "000000010111100011111101010" OR uut_a_5_5 /= "000000000010011010010110111" THEN
              FAIL <= '1';
              FAIL_NUM <= "10011100";
              state <= "11111101";
            ELSE
              state <= "10101010";
            END IF;
            uut_rst <= '0';
          WHEN "10101010" =>
            uut_coord_shift <= "0111";
            uut_x <= "111100001011";
            uut_y <= "111111011111";
            uut_fx <= "0101010100";
            uut_fy <= "0001111000";
            uut_ft <= "0000010101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000010011001111010100100" OR uut_a_0_1 /= "111111101100110000101011100" OR uut_a_0_2 /= "101111100111011101000010110" OR uut_a_0_3 /= "111111101010011000101101000" OR uut_a_0_4 /= "000000010101100111010011000" OR uut_a_0_5 /= "010010011001111101101011100" OR uut_a_1_0 /= "111111111111101100110000101" OR uut_a_1_1 /= "000000000000010011001111010" OR uut_a_1_2 /= "000000010000011000100010111" OR uut_a_1_3 /= "000000000000010101100111010" OR uut_a_1_4 /= "111111111111101010011000101" OR uut_a_1_5 /= "111111101101100110000010010" OR uut_a_2_0 /= "111111101111100111011101000" OR uut_a_2_1 /= "000000010000011000100010111" OR uut_a_2_2 /= "001101111100111001110001001" OR uut_a_2_3 /= "000000010010011001111101101" OR uut_a_2_4 /= "111111101101100110000010010" OR uut_a_2_5 /= "110000010100111000111110011" OR uut_a_3_0 /= "111111101010011000101101000" OR uut_a_3_1 /= "000000010101100111010011000" OR uut_a_3_2 /= "010010011001111101101011100" OR uut_a_3_3 /= "000000011000010010000010000" OR uut_a_3_4 /= "111111100111101101111110000" OR uut_a_3_5 /= "101011010100101001010011000" OR uut_a_4_0 /= "000000000000010101100111010" OR uut_a_4_1 /= "111111111111101010011000101" OR uut_a_4_2 /= "111111101101100110000010010" OR uut_a_4_3 /= "111111111111100111101101111" OR uut_a_4_4 /= "000000000000011000010010000" OR uut_a_4_5 /= "000000010100101011010110101" OR uut_a_5_0 /= "000000010010011001111101101" OR uut_a_5_1 /= "111111101101100110000010010" OR uut_a_5_2 /= "110000010100111000111110011" OR uut_a_5_3 /= "111111101011010100101001010" OR uut_a_5_4 /= "000000010100101011010110101" OR uut_a_5_5 /= "010001100110111010110101010" THEN
              FAIL <= '1';
              FAIL_NUM <= "10011101";
              state <= "11111101";
            ELSE
              state <= "10101011";
            END IF;
            uut_rst <= '0';
          WHEN "10101011" =>
            uut_coord_shift <= "0111";
            uut_x <= "000010111010";
            uut_y <= "111100110011";
            uut_fx <= "0110100010";
            uut_fy <= "1001101111";
            uut_ft <= "0000010001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001101001001000000" OR uut_a_0_1 /= "000001000100001010101100000" OR uut_a_0_2 /= "111111101010101001011000000" OR uut_a_0_3 /= "000000000100100111011100000" OR uut_a_0_4 /= "000010111111100100101010000" OR uut_a_0_5 /= "111111000011111111010100000" OR uut_a_1_0 /= "000000000001000100001010101" OR uut_a_1_1 /= "000000101100001100111011100" OR uut_a_1_2 /= "111111110010001001110101000" OR uut_a_1_3 /= "000000000010111111100100101" OR uut_a_1_4 /= "000001111100001110010001001" OR uut_a_1_5 /= "111111011001000101100011011" OR uut_a_2_0 /= "111111111111101010101001011" OR uut_a_2_1 /= "111111110010001001110101000" OR uut_a_2_2 /= "000000000100010101100110001" OR uut_a_2_3 /= "111111111111000011111111010" OR uut_a_2_4 /= "111111011001000101100011011" OR uut_a_2_5 /= "000000001100001100001000111" OR uut_a_3_0 /= "000000000100100111011100000" OR uut_a_3_1 /= "000010111111100100101010000" OR uut_a_3_2 /= "111111000011111111010100000" OR uut_a_3_3 /= "000000001100111110010010000" OR uut_a_3_4 /= "001000011010011000101011000" OR uut_a_3_5 /= "111101010111010110010110000" OR uut_a_4_0 /= "000000000010111111100100101" OR uut_a_4_1 /= "000001111100001110010001001" OR uut_a_4_2 /= "111111011001000101100011011" OR uut_a_4_3 /= "000000001000011010011000101" OR uut_a_4_4 /= "000101011101000110111111111" OR uut_a_4_5 /= "111110010010101000111111010" OR uut_a_5_0 /= "111111111111000011111111010" OR uut_a_5_1 /= "111111011001000101100011011" OR uut_a_5_2 /= "000000001100001100001000111" OR uut_a_5_3 /= "111111111101010111010110010" OR uut_a_5_4 /= "111110010010101000111111010" OR uut_a_5_5 /= "000000100010010000011101100" THEN
              FAIL <= '1';
              FAIL_NUM <= "10011110";
              state <= "11111101";
            ELSE
              state <= "10101100";
            END IF;
            uut_rst <= '0';
          WHEN "10101100" =>
            uut_coord_shift <= "0111";
            uut_x <= "111101001010";
            uut_y <= "000000011110";
            uut_fx <= "1000000101";
            uut_fy <= "0100010001";
            uut_ft <= "0101100101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000111011100101000100" OR uut_a_0_1 /= "000110011001100110110011100" OR uut_a_0_2 /= "111011011001110101000000010" OR uut_a_0_3 /= "111111110011101110100111100" OR uut_a_0_4 /= "110101011101000011111100100" OR uut_a_0_5 /= "000111100100101110100111110" OR uut_a_1_0 /= "000000000110011001100110110" OR uut_a_1_1 /= "000101100000000000010110010" OR uut_a_1_2 /= "111100000011001100100011001" OR uut_a_1_3 /= "111111110101011101000011111" OR uut_a_1_4 /= "110110111011111110011000111" OR uut_a_1_5 /= "000110100000100100000100001" OR uut_a_2_0 /= "111111111011011001110101000" OR uut_a_2_1 /= "111100000011001100100011001" OR uut_a_2_2 /= "000010110101100011110010010" OR uut_a_2_3 /= "000000000111100100101110100" OR uut_a_2_4 /= "000110100000100100000100001" OR uut_a_2_5 /= "111011010100110101001110011" OR uut_a_3_0 /= "111111110011101110100111100" OR uut_a_3_1 /= "110101011101000011111100100" OR uut_a_3_2 /= "000111100100101110100111110" OR uut_a_3_3 /= "000000010100001110001000100" OR uut_a_3_4 /= "010001011000001001010011100" OR uut_a_3_5 /= "110011100001010001110000010" OR uut_a_4_0 /= "111111110101011101000011111" OR uut_a_4_1 /= "110110111011111110011000111" OR uut_a_4_2 /= "000110100000100100000100001" OR uut_a_4_3 /= "000000010001011000001001010" OR uut_a_4_4 /= "001110111011101111111111110" OR uut_a_4_5 /= "110101010001100110010000011" OR uut_a_5_0 /= "000000000111100100101110100" OR uut_a_5_1 /= "000110100000100100000100001" OR uut_a_5_2 /= "111011010100110101001110011" OR uut_a_5_3 /= "111111110011100001010001110" OR uut_a_5_4 /= "110101010001100110010000011" OR uut_a_5_5 /= "000111101100111101100010101" THEN
              FAIL <= '1';
              FAIL_NUM <= "10011111";
              state <= "11111101";
            ELSE
              state <= "10101101";
            END IF;
            uut_rst <= '0';
          WHEN "10101101" =>
            uut_coord_shift <= "0111";
            uut_x <= "000011010101";
            uut_y <= "000011111001";
            uut_fx <= "0000000101";
            uut_fy <= "1100010110";
            uut_ft <= "1001100111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000110100001101100010" OR uut_a_0_1 /= "000000000011010000110110001" OR uut_a_0_2 /= "000010111010000000001101001" OR uut_a_0_3 /= "000000000000101010001001110" OR uut_a_0_4 /= "000000000000010101000100111" OR uut_a_0_5 /= "000000010010110001010101111" OR uut_a_1_0 /= "000000000000000001101000011" OR uut_a_1_1 /= "000000000000000000110100001" OR uut_a_1_2 /= "000000000000101110100000000" OR uut_a_1_3 /= "000000000000000000001010100" OR uut_a_1_4 /= "000000000000000000000101010" OR uut_a_1_5 /= "000000000000000100101100010" OR uut_a_2_0 /= "000000000001011101000000000" OR uut_a_2_1 /= "000000000000101110100000000" OR uut_a_2_2 /= "000000101001011010100010111" OR uut_a_2_3 /= "000000000000001001011000101" OR uut_a_2_4 /= "000000000000000100101100010" OR uut_a_2_5 /= "000000000100001011011111000" OR uut_a_3_0 /= "000000000000101010001001110" OR uut_a_3_1 /= "000000000000010101000100111" OR uut_a_3_2 /= "000000010010110001010101111" OR uut_a_3_3 /= "000000000000000100010000010" OR uut_a_3_4 /= "000000000000000010001000001" OR uut_a_3_5 /= "000000000001111001001111001" OR uut_a_4_0 /= "000000000000000000001010100" OR uut_a_4_1 /= "000000000000000000000101010" OR uut_a_4_2 /= "000000000000000100101100010" OR uut_a_4_3 /= "000000000000000000000001000" OR uut_a_4_4 /= "000000000000000000000000100" OR uut_a_4_5 /= "000000000000000000011110010" OR uut_a_5_0 /= "000000000000001001011000101" OR uut_a_5_1 /= "000000000000000100101100010" OR uut_a_5_2 /= "000000000100001011011111000" OR uut_a_5_3 /= "000000000000000000111100100" OR uut_a_5_4 /= "000000000000000000011110010" OR uut_a_5_5 /= "000000000000011010111111100" THEN
              FAIL <= '1';
              FAIL_NUM <= "10100000";
              state <= "11111101";
            ELSE
              state <= "10101110";
            END IF;
            uut_rst <= '0';
          WHEN "10101110" =>
            uut_coord_shift <= "0111";
            uut_x <= "000000000100";
            uut_y <= "000000101011";
            uut_fx <= "0100001101";
            uut_fy <= "1001010101";
            uut_ft <= "0010100101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000001101111000110010010" OR uut_a_0_1 /= "111101100000010010111110001" OR uut_a_0_2 /= "111100000110000001110111100" OR uut_a_0_3 /= "000000000011100101001011110" OR uut_a_0_4 /= "111111010110110100011000111" OR uut_a_0_5 /= "111110111111100010101100100" OR uut_a_1_0 /= "111111111110110000001001011" OR uut_a_1_1 /= "000000001110010110010010111" OR uut_a_1_2 /= "000000010110011101010101010" OR uut_a_1_3 /= "111111111111101011011010001" OR uut_a_1_4 /= "000000000011101100110010110" OR uut_a_1_5 /= "000000000101110010101000100" OR uut_a_2_0 /= "111111111110000011000000111" OR uut_a_2_1 /= "000000010110011101010101010" OR uut_a_2_2 /= "000000100011001001101111001" OR uut_a_2_3 /= "111111111111011111110001010" OR uut_a_2_4 /= "000000000101110010101000100" OR uut_a_2_5 /= "000000001001000100000111101" OR uut_a_3_0 /= "000000000011100101001011110" OR uut_a_3_1 /= "111111010110110100011000111" OR uut_a_3_2 /= "111110111111100010101100100" OR uut_a_3_3 /= "000000000000111011000110010" OR uut_a_3_4 /= "111111110101011000011000001" OR uut_a_3_5 /= "111111101111011000001111100" OR uut_a_4_0 /= "111111111111101011011010001" OR uut_a_4_1 /= "000000000011101100110010110" OR uut_a_4_2 /= "000000000101110010101000100" OR uut_a_4_3 /= "111111111111111010101100001" OR uut_a_4_4 /= "000000000000111101000011110" OR uut_a_4_5 /= "000000000001011111100100100" OR uut_a_5_0 /= "111111111111011111110001010" OR uut_a_5_1 /= "000000000101110010101000100" OR uut_a_5_2 /= "000000001001000100000111101" OR uut_a_5_3 /= "111111111111110111101100000" OR uut_a_5_4 /= "000000000001011111100100100" OR uut_a_5_5 /= "000000000010010101100101110" THEN
              FAIL <= '1';
              FAIL_NUM <= "10100001";
              state <= "11111101";
            ELSE
              state <= "10101111";
            END IF;
            uut_rst <= '0';
          WHEN "10101111" =>
            uut_coord_shift <= "0111";
            uut_x <= "000000001000";
            uut_y <= "111101011000";
            uut_fx <= "0111000001";
            uut_fy <= "0001011101";
            uut_ft <= "1111000011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000001001000010" OR uut_a_0_1 /= "000000000000111111001110000" OR uut_a_0_2 /= "111111111111010011111110010" OR uut_a_0_3 /= "000000000000000011110110100" OR uut_a_0_4 /= "000000000011010111101100000" OR uut_a_0_5 /= "111111111101101001110010100" OR uut_a_1_0 /= "000000000000000000011111100" OR uut_a_1_1 /= "000000000000011011101010001" OR uut_a_1_2 /= "111111111111101100101111001" OR uut_a_1_3 /= "000000000000000001101011110" OR uut_a_1_4 /= "000000000001011110010111010" OR uut_a_1_5 /= "111111111110111110010010000" OR uut_a_2_0 /= "111111111111111111101001111" OR uut_a_2_1 /= "111111111111101100101111001" OR uut_a_2_2 /= "000000000000001101011010100" OR uut_a_2_3 /= "111111111111111110110100111" OR uut_a_2_4 /= "111111111110111110010010000" OR uut_a_2_5 /= "000000000000101101110001000" OR uut_a_3_0 /= "000000000000000011110110100" OR uut_a_3_1 /= "000000000011010111101100000" OR uut_a_3_2 /= "111111111101101001110010100" OR uut_a_3_3 /= "000000000000001101001001000" OR uut_a_3_4 /= "000000001011011111111000000" OR uut_a_3_5 /= "111111110111111111100001000" OR uut_a_4_0 /= "000000000000000001101011110" OR uut_a_4_1 /= "000000000001011110010111010" OR uut_a_4_2 /= "111111111110111110010010000" OR uut_a_4_3 /= "000000000000000101101111111" OR uut_a_4_4 /= "000000000101000001111100100" OR uut_a_4_5 /= "111111111100011111110010011" OR uut_a_5_0 /= "111111111111111110110100111" OR uut_a_5_1 /= "111111111110111110010010000" OR uut_a_5_2 /= "000000000000101101110001000" OR uut_a_5_3 /= "111111111111111011111111110" OR uut_a_5_4 /= "111111111100011111110010011" OR uut_a_5_5 /= "000000000010011100001001011" THEN
              FAIL <= '1';
              FAIL_NUM <= "10100010";
              state <= "11111101";
            ELSE
              state <= "10110000";
            END IF;
            uut_rst <= '0';
          WHEN "10110000" =>
            uut_coord_shift <= "0111";
            uut_x <= "000011100010";
            uut_y <= "000001001111";
            uut_fx <= "1111001111";
            uut_fy <= "0101011100";
            uut_ft <= "0000100001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000010101111110010" OR uut_a_0_1 /= "000000000101010100100100111" OR uut_a_0_2 /= "000000010000111111101001011" OR uut_a_0_3 /= "111111111110011011001110000" OR uut_a_0_4 /= "111111100111100101111001000" OR uut_a_0_5 /= "111110110010000011010101000" OR uut_a_1_0 /= "000000000000000010101010010" OR uut_a_1_1 /= "000000000000101001001111011" OR uut_a_1_2 /= "000000000010000011101101010" OR uut_a_1_3 /= "111111111111110011110010111" OR uut_a_1_4 /= "111111111101000010110101101" OR uut_a_1_5 /= "111111110110100011111001110" OR uut_a_2_0 /= "000000000000001000011111110" OR uut_a_2_1 /= "000000000010000011101101010" OR uut_a_2_2 /= "000000000110100100100111010" OR uut_a_2_3 /= "111111111111011001000001101" OR uut_a_2_4 /= "111111110110100011111001110" OR uut_a_2_5 /= "111111100001110110110010010" OR uut_a_3_0 /= "111111111110011011001110000" OR uut_a_3_1 /= "111111100111100101111001000" OR uut_a_3_2 /= "111110110010000011010101000" OR uut_a_3_3 /= "000000000111001110010000000" OR uut_a_3_4 /= "000001101111111100111000000" OR uut_a_3_5 /= "000101100101100001011000000" OR uut_a_4_0 /= "111111111111110011110010111" OR uut_a_4_1 /= "111111111101000010110101101" OR uut_a_4_2 /= "111111110110100011111001110" OR uut_a_4_3 /= "000000000000110111111110011" OR uut_a_4_4 /= "000000001101100011100111110" OR uut_a_4_5 /= "000000101011010010110010101" OR uut_a_5_0 /= "111111111111011001000001101" OR uut_a_5_1 /= "111111110110100011111001110" OR uut_a_5_2 /= "111111100001110110110010010" OR uut_a_5_3 /= "000000000010110010110000101" OR uut_a_5_4 /= "000000101011010010110010101" OR uut_a_5_5 /= "000010001010010000101010000" THEN
              FAIL <= '1';
              FAIL_NUM <= "10100011";
              state <= "11111101";
            ELSE
              state <= "10110001";
            END IF;
            uut_rst <= '0';
          WHEN "10110001" =>
            uut_coord_shift <= "0111";
            uut_x <= "000000011011";
            uut_y <= "000001011100";
            uut_fx <= "1101111000";
            uut_fy <= "1011110101";
            uut_ft <= "0001010001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000110100100100000" OR uut_a_0_1 /= "111111100010110110000010000" OR uut_a_0_2 /= "111111110110100011100010000" OR uut_a_0_3 /= "111111111110000000001110000" OR uut_a_0_4 /= "000001000110111000001111000" OR uut_a_0_5 /= "000000010110111101011111000" OR uut_a_1_0 /= "111111111111110001011011000" OR uut_a_1_1 /= "000000001000000101100000111" OR uut_a_1_2 /= "000000000010100111101001010" OR uut_a_1_3 /= "000000000000100011011100000" OR uut_a_1_4 /= "111111101100010101111001110" OR uut_a_1_5 /= "111111111001101000011100101" OR uut_a_2_0 /= "111111111111111011010001110" OR uut_a_2_1 /= "000000000010100111101001010" OR uut_a_2_2 /= "000000000000110110010011101" OR uut_a_2_3 /= "000000000000001011011110101" OR uut_a_2_4 /= "111111111001101000011100101" OR uut_a_2_5 /= "111111111101111011111110011" OR uut_a_3_0 /= "111111111110000000001110000" OR uut_a_3_1 /= "000001000110111000001111000" OR uut_a_3_2 /= "000000010110111101011111000" OR uut_a_3_3 /= "000000000100110110101001000" OR uut_a_3_4 /= "111101010011101100010000100" OR uut_a_3_5 /= "111111001000001011101000100" OR uut_a_4_0 /= "000000000000100011011100000" OR uut_a_4_1 /= "111111101100010101111001110" OR uut_a_4_2 /= "111111111001101000011100101" OR uut_a_4_3 /= "111111111110101001110110001" OR uut_a_4_4 /= "000000101111110010011110011" OR uut_a_4_5 /= "000000001111011110110001100" OR uut_a_5_0 /= "000000000000001011011110101" OR uut_a_5_1 /= "111111111001101000011100101" OR uut_a_5_2 /= "111111111101111011111110011" OR uut_a_5_3 /= "111111111111100100000101110" OR uut_a_5_4 /= "000000001111011110110001100" OR uut_a_5_5 /= "000000000101000000111101000" THEN
              FAIL <= '1';
              FAIL_NUM <= "10100100";
              state <= "11111101";
            ELSE
              state <= "10110010";
            END IF;
            uut_rst <= '0';
          WHEN "10110010" =>
            uut_coord_shift <= "0111";
            uut_x <= "000010111011";
            uut_y <= "111111010001";
            uut_fx <= "1001110011";
            uut_fy <= "1111000110";
            uut_ft <= "1100110011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000001100101100010000000" OR uut_a_0_1 /= "111100100001111001101000000" OR uut_a_0_2 /= "001001110100001110011000000" OR uut_a_0_3 /= "000000001000000110010110000" OR uut_a_0_4 /= "111101110010010000111111000" OR uut_a_0_5 /= "000110010000111010000001000" OR uut_a_1_0 /= "111111111110010000111100110" OR uut_a_1_1 /= "000000011110010111010111110" OR uut_a_1_2 /= "111110101010000111000010001" OR uut_a_1_3 /= "111111111110111001001000011" OR uut_a_1_4 /= "000000010011011000001011011" OR uut_a_1_5 /= "111111001001001100000100010" OR uut_a_2_0 /= "000000000100111010000111001" OR uut_a_2_1 /= "111110101010000111000010001" OR uut_a_2_2 /= "000011110010111100100011110" OR uut_a_2_3 /= "000000000011001000011101000" OR uut_a_2_4 /= "111111001001001100000100010" OR uut_a_2_5 /= "000010011011000010011011111" OR uut_a_3_0 /= "000000001000000110010110000" OR uut_a_3_1 /= "111101110010010000111111000" OR uut_a_3_2 /= "000110010000111010000001000" OR uut_a_3_3 /= "000000000101001010110010010" OR uut_a_3_4 /= "111110100101100011010000101" OR uut_a_3_5 /= "000011111111110101110111011" OR uut_a_4_0 /= "111111111110111001001000011" OR uut_a_4_1 /= "000000010011011000001011011" OR uut_a_4_2 /= "111111001001001100000100010" OR uut_a_4_3 /= "111111111111010010110001101" OR uut_a_4_4 /= "000000001100010111011011011" OR uut_a_4_5 /= "111111011101000001011000101" OR uut_a_5_0 /= "000000000011001000011101000" OR uut_a_5_1 /= "111111001001001100000100010" OR uut_a_5_2 /= "000010011011000010011011111" OR uut_a_5_3 /= "000000000001111111111010111" OR uut_a_5_4 /= "111111011101000001011000101" OR uut_a_5_5 /= "000001100010111100000101001" THEN
              FAIL <= '1';
              FAIL_NUM <= "10100101";
              state <= "11111101";
            ELSE
              state <= "10110011";
            END IF;
            uut_rst <= '0';
          WHEN "10110011" =>
            uut_coord_shift <= "0111";
            uut_x <= "111111001110";
            uut_y <= "000010101010";
            uut_fx <= "1110011101";
            uut_fy <= "1110010000";
            uut_ft <= "1101110001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000100001110010010" OR uut_a_0_1 /= "111111001011001101011111000" OR uut_a_0_2 /= "111111110001001110000001000" OR uut_a_0_3 /= "111111111111110000101111100" OR uut_a_0_4 /= "000000010111110101110010000" OR uut_a_0_5 /= "000000000110101011001110000" OR uut_a_1_0 /= "111111111111100101100110101" OR uut_a_1_1 /= "000000101001001111011101110" OR uut_a_1_2 /= "000000001011100011000011001" OR uut_a_1_3 /= "000000000000001011111010111" OR uut_a_1_4 /= "111111101101010111111110111" OR uut_a_1_5 /= "111111111010110010001111000" OR uut_a_2_0 /= "111111111111111000100111000" OR uut_a_2_1 /= "000000001011100011000011001" OR uut_a_2_2 /= "000000000011001110111011110" OR uut_a_2_3 /= "000000000000000011010101100" OR uut_a_2_4 /= "111111111010110010001111000" OR uut_a_2_5 /= "111111111110100010100010111" OR uut_a_3_0 /= "111111111111110000101111100" OR uut_a_3_1 /= "000000010111110101110010000" OR uut_a_3_2 /= "000000000110101011001110000" OR uut_a_3_3 /= "000000000000000110111001000" OR uut_a_3_4 /= "111111110101001110111100000" OR uut_a_3_5 /= "111111111100111111000100000" OR uut_a_4_0 /= "000000000000001011111010111" OR uut_a_4_1 /= "111111101101010111111110111" OR uut_a_4_2 /= "111111111010110010001111000" OR uut_a_4_3 /= "111111111111111010100111011" OR uut_a_4_4 /= "000000001000011010010101001" OR uut_a_4_5 /= "000000000010010110101110111" OR uut_a_5_0 /= "000000000000000011010101100" OR uut_a_5_1 /= "111111111010110010001111000" OR uut_a_5_2 /= "111111111110100010100010111" OR uut_a_5_3 /= "111111111111111110011111100" OR uut_a_5_4 /= "000000000010010110101110111" OR uut_a_5_5 /= "000000000000101010001101001" THEN
              FAIL <= '1';
              FAIL_NUM <= "10100110";
              state <= "11111101";
            ELSE
              state <= "10110100";
            END IF;
            uut_rst <= '0';
          WHEN "10110100" =>
            uut_coord_shift <= "1000";
            uut_x <= "111010010000";
            uut_y <= "111100001011";
            uut_fx <= "1001011001";
            uut_fy <= "1110111000";
            uut_ft <= "1100000111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000001111000001000000000" OR uut_a_0_1 /= "101111110011111011000000000" OR uut_a_0_2 /= "010100000011110101100000000" OR uut_a_0_3 /= "111111110100101111010000000" OR uut_a_0_4 /= "001100001001000011110000000" OR uut_a_0_5 /= "110000111101000111111000000" OR uut_a_1_0 /= "111111110111111001111101100" OR uut_a_1_1 /= "001000101110100000101100100" OR uut_a_1_2 /= "110101001011111011101010010" OR uut_a_1_3 /= "000000000110000100100001111" OR uut_a_1_4 /= "111001011101000111011110101" OR uut_a_1_5 /= "001000000111000011010000010" OR uut_a_2_0 /= "000000001010000001111010110" OR uut_a_2_1 /= "110101001011111011101010010" OR uut_a_2_2 /= "001101011001100011111111001" OR uut_a_2_3 /= "111111111000011110100011111" OR uut_a_2_4 /= "001000000111000011010000010" OR uut_a_2_5 /= "110101111100110101000000101" OR uut_a_3_0 /= "111111110100101111010000000" OR uut_a_3_1 /= "001100001001000011110000000" OR uut_a_3_2 /= "110000111101000111111000000" OR uut_a_3_3 /= "000000001000011100100100000" OR uut_a_3_4 /= "110110111001001101001100000" OR uut_a_3_5 /= "001011010010001010000110000" OR uut_a_4_0 /= "000000000110000100100001111" OR uut_a_4_1 /= "111001011101000111011110101" OR uut_a_4_2 /= "001000000111000011010000010" OR uut_a_4_3 /= "111111111011011100100110100" OR uut_a_4_4 /= "000100111010001010011001000" OR uut_a_4_5 /= "111001111010101101100011110" OR uut_a_5_0 /= "111111111000011110100011111" OR uut_a_5_1 /= "001000000111000011010000010" OR uut_a_5_2 /= "110101111100110101000000101" OR uut_a_5_3 /= "000000000101101001000101000" OR uut_a_5_4 /= "111001111010101101100011110" OR uut_a_5_5 /= "000111100010011000001111100" THEN
              FAIL <= '1';
              FAIL_NUM <= "10100111";
              state <= "11111101";
            ELSE
              state <= "10110101";
            END IF;
            uut_rst <= '0';
          WHEN "10110101" =>
            uut_coord_shift <= "1000";
            uut_x <= "111100110001";
            uut_y <= "111110110100";
            uut_fx <= "1001111010";
            uut_fy <= "1111111011";
            uut_ft <= "0011010011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000101000110010000010" OR uut_a_0_1 /= "000011011011001100111010110" OR uut_a_0_2 /= "000000000000000000000000000" OR uut_a_0_3 /= "111111111110101101100101110" OR uut_a_0_4 /= "111111001000101000010111010" OR uut_a_0_5 /= "000000000000000000000000000" OR uut_a_1_0 /= "000000000001101101100110011" OR uut_a_1_1 /= "000001001001101000110101101" OR uut_a_1_2 /= "000000000000000000000000000" OR uut_a_1_3 /= "111111111111100100010100001" OR uut_a_1_4 /= "111111101101011001100011110" OR uut_a_1_5 /= "000000000000000000000000000" OR uut_a_2_0 /= "000000000000000000000000000" OR uut_a_2_1 /= "000000000000000000000000000" OR uut_a_2_2 /= "000000000000000000000000000" OR uut_a_2_3 /= "000000000000000000000000000" OR uut_a_2_4 /= "000000000000000000000000000" OR uut_a_2_5 /= "000000000000000000000000000" OR uut_a_3_0 /= "111111111110101101100101110" OR uut_a_3_1 /= "111111001000101000010111010" OR uut_a_3_2 /= "000000000000000000000000000" OR uut_a_3_3 /= "000000000000010100110100010" OR uut_a_3_4 /= "000000001101111111000110110" OR uut_a_3_5 /= "000000000000000000000000000" OR uut_a_4_0 /= "111111111111100100010100001" OR uut_a_4_1 /= "111111101101011001100011110" OR uut_a_4_2 /= "000000000000000000000000000" OR uut_a_4_3 /= "000000000000000110111111100" OR uut_a_4_4 /= "000000000100101100101100110" OR uut_a_4_5 /= "000000000000000000000000000" OR uut_a_5_0 /= "000000000000000000000000000" OR uut_a_5_1 /= "000000000000000000000000000" OR uut_a_5_2 /= "000000000000000000000000000" OR uut_a_5_3 /= "000000000000000000000000000" OR uut_a_5_4 /= "000000000000000000000000000" OR uut_a_5_5 /= "000000000000000000000000000" THEN
              FAIL <= '1';
              FAIL_NUM <= "10101000";
              state <= "11111101";
            ELSE
              state <= "10110110";
            END IF;
            uut_rst <= '0';
          WHEN "10110110" =>
            uut_coord_shift <= "1000";
            uut_x <= "111011111010";
            uut_y <= "000100100011";
            uut_fx <= "1001001100";
            uut_fy <= "1110010011";
            uut_ft <= "1000000011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000001100101000101100010" OR uut_a_0_1 /= "001000100101101010000100111" OR uut_a_0_2 /= "000100111011111001010010010" OR uut_a_0_3 /= "000000001100100110111010100" OR uut_a_0_4 /= "001000100100011100110000110" OR uut_a_0_5 /= "000100111011001100110110100" OR uut_a_1_0 /= "000000000100010010110101000" OR uut_a_1_1 /= "000010111010110011000011001" OR uut_a_1_2 /= "000001101011010110101101111" OR uut_a_1_3 /= "000000000100010010001110011" OR uut_a_1_4 /= "000010111010011000110001100" OR uut_a_1_5 /= "000001101011000111100111100" OR uut_a_2_0 /= "000000000010011101111100101" OR uut_a_2_1 /= "000001101011010110101101111" OR uut_a_2_2 /= "000000111101101100101100000" OR uut_a_2_3 /= "000000000010011101100110011" OR uut_a_2_4 /= "000001101011000111100111100" OR uut_a_2_5 /= "000000111101100100000000101" OR uut_a_3_0 /= "000000001100100110111010100" OR uut_a_3_1 /= "001000100100011100110000110" OR uut_a_3_2 /= "000100111011001100110110100" OR uut_a_3_3 /= "000000001100100101001001000" OR uut_a_3_4 /= "001000100011001111100111100" OR uut_a_3_5 /= "000100111010100000100001000" OR uut_a_4_0 /= "000000000100010010001110011" OR uut_a_4_1 /= "000010111010011000110001100" OR uut_a_4_2 /= "000001101011000111100111100" OR uut_a_4_3 /= "000000000100010001100111110" OR uut_a_4_4 /= "000010111001111110100011101" OR uut_a_4_5 /= "000001101010111000100011001" OR uut_a_5_0 /= "000000000010011101100110011" OR uut_a_5_1 /= "000001101011000111100111100" OR uut_a_5_2 /= "000000111101100100000000101" OR uut_a_5_3 /= "000000000010011101010000010" OR uut_a_5_4 /= "000001101010111000100011001" OR uut_a_5_5 /= "000000111101011011010110011" THEN
              FAIL <= '1';
              FAIL_NUM <= "10101001";
              state <= "11111101";
            ELSE
              state <= "10110111";
            END IF;
            uut_rst <= '0';
          WHEN "10110111" =>
            uut_coord_shift <= "1000";
            uut_x <= "111011100010";
            uut_y <= "111000000010";
            uut_fx <= "1011000010";
            uut_fy <= "1010010010";
            uut_ft <= "1100010011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000111000011100100000" OR uut_a_0_1 /= "110010011111101011100110000" OR uut_a_0_2 /= "111110001011100101001110000" OR uut_a_0_3 /= "000000000010011111011000000" OR uut_a_0_4 /= "111011001110111100100100000" OR uut_a_0_5 /= "111111010110111010010100000" OR uut_a_1_0 /= "111111111001001111110101110" OR uut_a_1_1 /= "001100111011001011100001111" OR uut_a_1_2 /= "000001101111011010101000010" OR uut_a_1_3 /= "111111111101100111011110010" OR uut_a_1_4 /= "000100100011111100100010100" OR uut_a_1_5 /= "000000100111010100101100010" OR uut_a_2_0 /= "111111111111000101110010100" OR uut_a_2_1 /= "000001101111011010101000010" OR uut_a_2_2 /= "000000001111000000011100111" OR uut_a_2_3 /= "111111111111101011011101001" OR uut_a_2_4 /= "000000100111010100101100010" OR uut_a_2_5 /= "000000000101010010111110111" OR uut_a_3_0 /= "000000000010011111011000000" OR uut_a_3_1 /= "111011001110111100100100000" OR uut_a_3_2 /= "111111010110111010010100000" OR uut_a_3_3 /= "000000000000111000010000000" OR uut_a_3_4 /= "111110010100010101011000000" OR uut_a_3_5 /= "111111110001011111111000000" OR uut_a_4_0 /= "111111111101100111011110010" OR uut_a_4_1 /= "000100100011111100100010100" OR uut_a_4_2 /= "000000100111010100101100010" OR uut_a_4_3 /= "111111111111001010001010101" OR uut_a_4_4 /= "000001100111000010100010110" OR uut_a_4_5 /= "000000001101111000001111101" OR uut_a_5_0 /= "111111111111101011011101001" OR uut_a_5_1 /= "000000100111010100101100010" OR uut_a_5_2 /= "000000000101010010111110111" OR uut_a_5_3 /= "111111111111111000101111111" OR uut_a_5_4 /= "000000001101111000001111101" OR uut_a_5_5 /= "000000000001110111101001000" THEN
              FAIL <= '1';
              FAIL_NUM <= "10101010";
              state <= "11111101";
            ELSE
              state <= "10111000";
            END IF;
            uut_rst <= '0';
          WHEN "10111000" =>
            uut_coord_shift <= "1000";
            uut_x <= "111010110100";
            uut_y <= "111010001110";
            uut_fx <= "0001100101";
            uut_fy <= "0110011011";
            uut_ft <= "0111000010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000001010101010100001000" OR uut_a_0_1 /= "001111011111110001111101000" OR uut_a_0_2 /= "101110111010111010001001100" OR uut_a_0_3 /= "111111110101110001001111100" OR uut_a_0_4 /= "110001001000100011100001100" OR uut_a_0_5 /= "010000011000101000101011010" OR uut_a_1_0 /= "000000000111101111111000111" OR uut_a_1_1 /= "001011010000100101110010110" OR uut_a_1_2 /= "110011100101110011001111111" OR uut_a_1_3 /= "111111111000100100010001110" OR uut_a_1_4 /= "110101001100101101110011110" OR uut_a_1_5 /= "001011111001111001100011011" OR uut_a_2_0 /= "111111110111011101011101000" OR uut_a_2_1 /= "110011100101110011001111111" OR uut_a_2_2 /= "001101101011010100111011111" OR uut_a_2_3 /= "000000001000001100010100010" OR uut_a_2_4 /= "001011111001111001100011011" OR uut_a_2_5 /= "110010111000010001011011010" OR uut_a_3_0 /= "111111110101110001001111100" OR uut_a_3_1 /= "110001001000100011100001100" OR uut_a_3_2 /= "010000011000101000101011010" OR uut_a_3_3 /= "000000001001110100001000010" OR uut_a_3_4 /= "001110010000101111111111010" OR uut_a_3_5 /= "110000010010000000110010011" OR uut_a_4_0 /= "111111111000100100010001110" OR uut_a_4_1 /= "110101001100101101110011110" OR uut_a_4_2 /= "001011111001111001100011011" OR uut_a_4_3 /= "000000000111001000010111111" OR uut_a_4_4 /= "001010010111001010110111011" OR uut_a_4_5 /= "110100100101000101100100100" OR uut_a_5_0 /= "000000001000001100010100010" OR uut_a_5_1 /= "001011111001111001100011011" OR uut_a_5_2 /= "110010111000010001011011010" OR uut_a_5_3 /= "111111111000001001000000011" OR uut_a_5_4 /= "110100100101000101100100100" OR uut_a_5_5 /= "001100100101100100110111101" THEN
              FAIL <= '1';
              FAIL_NUM <= "10101011";
              state <= "11111101";
            ELSE
              state <= "10111001";
            END IF;
            uut_rst <= '0';
          WHEN "10111001" =>
            uut_coord_shift <= "1000";
            uut_x <= "111011100011";
            uut_y <= "111111101111";
            uut_fx <= "1110000001";
            uut_fy <= "0000011000";
            uut_ft <= "1100001111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000001111101100000110010" OR uut_a_0_1 /= "101001101100010011000111010" OR uut_a_0_2 /= "000011101011010101011101110" OR uut_a_0_3 /= "111111110111100011010101010" OR uut_a_0_4 /= "001100000000110000110010010" OR uut_a_0_5 /= "111110000001010001111110110" OR uut_a_1_0 /= "111111110100110110001001100" OR uut_a_1_1 /= "001111110111000000011010010" OR uut_a_1_2 /= "111101011000101100001111010" OR uut_a_1_3 /= "000000000110000000011000011" OR uut_a_1_4 /= "110111011101011101010100010" OR uut_a_1_5 /= "000001011010000101101101111" OR uut_a_2_0 /= "000000000001110101101010101" OR uut_a_2_1 /= "111101011000101100001111010" OR uut_a_2_2 /= "000000011011100101000000111" OR uut_a_2_3 /= "111111111111000000101000111" OR uut_a_2_4 /= "000001011010000101101101111" OR uut_a_2_5 /= "111111110001001001100110110" OR uut_a_3_0 /= "111111110111100011010101010" OR uut_a_3_1 /= "001100000000110000110010010" OR uut_a_3_2 /= "111110000001010001111110110" OR uut_a_3_3 /= "000000000100100011001000010" OR uut_a_3_4 /= "111001100010000011010001010" OR uut_a_3_5 /= "000001000100001110111011110" OR uut_a_4_0 /= "000000000110000000011000011" OR uut_a_4_1 /= "110111011101011101010100010" OR uut_a_4_2 /= "000001011010000101101101111" OR uut_a_4_3 /= "111111111100110001000001101" OR uut_a_4_4 /= "000100100110010010101011001" OR uut_a_4_5 /= "111111001111011111011000100" OR uut_a_5_0 /= "111111111111000000101000111" OR uut_a_5_1 /= "000001011010000101101101111" OR uut_a_5_2 /= "111111110001001001100110110" OR uut_a_5_3 /= "000000000000100010000111011" OR uut_a_5_4 /= "111111001111011111011000100" OR uut_a_5_5 /= "000000000111111111110000000" THEN
              FAIL <= '1';
              FAIL_NUM <= "10101100";
              state <= "11111101";
            ELSE
              state <= "10111010";
            END IF;
            uut_rst <= '0';
          WHEN "10111010" =>
            uut_coord_shift <= "1000";
            uut_x <= "111001000110";
            uut_y <= "111110111111";
            uut_fx <= "1010110010";
            uut_fy <= "1000011011";
            uut_ft <= "0111010010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000000000110010" OR uut_a_0_1 /= "000000000000001010011001101" OR uut_a_0_2 /= "000000000000001100001010001" OR uut_a_0_3 /= "111111111111111011011011100" OR uut_a_0_4 /= "111111111000011001010000110" OR uut_a_0_5 /= "111111110111000110111111110" OR uut_a_1_0 /= "000000000000000000000101001" OR uut_a_1_1 /= "000000000000001000101001110" OR uut_a_1_2 /= "000000000000001010000111011" OR uut_a_1_3 /= "111111111111111100001100101" OR uut_a_1_4 /= "111111111001101011000001001" OR uut_a_1_5 /= "111111111000100110100100100" OR uut_a_2_0 /= "000000000000000000000110000" OR uut_a_2_1 /= "000000000000001010000111011" OR uut_a_2_2 /= "000000000000001011110100110" OR uut_a_2_3 /= "111111111111111011100011011" OR uut_a_2_4 /= "111111111000100110100100100" OR uut_a_2_5 /= "111111110111010110100011100" OR uut_a_3_0 /= "111111111111111011011011100" OR uut_a_3_1 /= "111111111000011001010000110" OR uut_a_3_2 /= "111111110111000110111111110" OR uut_a_3_3 /= "000000000011010101111001000" OR uut_a_3_4 /= "000101100011111011010110100" OR uut_a_3_5 /= "000110100000000101011000100" OR uut_a_4_0 /= "111111111111111100001100101" OR uut_a_4_1 /= "111111111001101011000001001" OR uut_a_4_2 /= "111111111000100110100100100" OR uut_a_4_3 /= "000000000010110001111101101" OR uut_a_4_4 /= "000100101000001001001000011" OR uut_a_4_5 /= "000101011010001100011110101" OR uut_a_5_0 /= "111111111111111011100011011" OR uut_a_5_1 /= "111111111000100110100100100" OR uut_a_5_2 /= "111111110111010110100011100" OR uut_a_5_3 /= "000000000011010000000010101" OR uut_a_5_4 /= "000101011010001100011110101" OR uut_a_5_5 /= "000110010100101101001111000" THEN
              FAIL <= '1';
              FAIL_NUM <= "10101101";
              state <= "11111101";
            ELSE
              state <= "10111011";
            END IF;
            uut_rst <= '0';
          WHEN "10111011" =>
            uut_coord_shift <= "1000";
            uut_x <= "111110111001";
            uut_y <= "000111011000";
            uut_fx <= "0100001101";
            uut_fy <= "1000001000";
            uut_ft <= "0010111000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000100011010101010010" OR uut_a_0_1 /= "000000001000110101010100100" OR uut_a_0_2 /= "000001011110111101001100011" OR uut_a_0_3 /= "111111111000111111010100010" OR uut_a_0_4 /= "111111110001111110101000100" OR uut_a_0_5 /= "111101101001010001010011011" OR uut_a_1_0 /= "000000000000000100011010101" OR uut_a_1_1 /= "000000000000001000110101010" OR uut_a_1_2 /= "000000000001011110111101001" OR uut_a_1_3 /= "111111111111111000111111010" OR uut_a_1_4 /= "111111111111110001111110101" OR uut_a_1_5 /= "111111111101101001010001010" OR uut_a_2_0 /= "000000000000101111011110100" OR uut_a_2_1 /= "000000000001011110111101001" OR uut_a_2_2 /= "000000001111111100110001110" OR uut_a_2_3 /= "111111111110110100101000101" OR uut_a_2_4 /= "111111111101101001010001010" OR uut_a_2_5 /= "111111100110101011101010000" OR uut_a_3_0 /= "111111111000111111010100010" OR uut_a_3_1 /= "111111110001111110101000100" OR uut_a_3_2 /= "111101101001010001010011011" OR uut_a_3_3 /= "000000001011001000001110010" OR uut_a_3_4 /= "000000010110010000011100100" OR uut_a_3_5 /= "000011101111010000110010011" OR uut_a_4_0 /= "111111111111111000111111010" OR uut_a_4_1 /= "111111111111110001111110101" OR uut_a_4_2 /= "111111111101101001010001010" OR uut_a_4_3 /= "000000000000001011001000001" OR uut_a_4_4 /= "000000000000010110010000011" OR uut_a_4_5 /= "000000000011101111010000110" OR uut_a_5_0 /= "111111111110110100101000101" OR uut_a_5_1 /= "111111111101101001010001010" OR uut_a_5_2 /= "111111100110101011101010000" OR uut_a_5_3 /= "000000000001110111101000011" OR uut_a_5_4 /= "000000000011101111010000110" OR uut_a_5_5 /= "000000101000001100000100011" THEN
              FAIL <= '1';
              FAIL_NUM <= "10101110";
              state <= "11111101";
            ELSE
              state <= "10111100";
            END IF;
            uut_rst <= '0';
          WHEN "10111100" =>
            uut_coord_shift <= "1000";
            uut_x <= "000011010010";
            uut_y <= "000010010100";
            uut_fx <= "0000110110";
            uut_fy <= "1011011111";
            uut_ft <= "0100010111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000001100010011100000010" OR uut_a_0_1 /= "000000110001001110000001000" OR uut_a_0_2 /= "101111110110011001101011000" OR uut_a_0_3 /= "000000000010100011000111010" OR uut_a_0_4 /= "000000001010001100011101000" OR uut_a_0_5 /= "111100101001111010011111000" OR uut_a_1_0 /= "000000000000011000100111000" OR uut_a_1_1 /= "000000000001100010011100000" OR uut_a_1_2 /= "111111011111101100110011010" OR uut_a_1_3 /= "000000000000000101000110001" OR uut_a_1_4 /= "000000000000010100011000111" OR uut_a_1_5 /= "111111111001010011110100111" OR uut_a_2_0 /= "111111110111111011001100110" OR uut_a_2_1 /= "111111011111101100110011010" OR uut_a_2_2 /= "001010100110010011001001110" OR uut_a_2_3 /= "111111111110010100111101001" OR uut_a_2_4 /= "111111111001010011110100111" OR uut_a_2_5 /= "000010001100011111100111101" OR uut_a_3_0 /= "000000000010100011000111010" OR uut_a_3_1 /= "000000001010001100011101000" OR uut_a_3_2 /= "111100101001111010011111000" OR uut_a_3_3 /= "000000000000100001110010010" OR uut_a_3_4 /= "000000000010000111001001000" OR uut_a_3_5 /= "111111010011101010000011000" OR uut_a_4_0 /= "000000000000000101000110001" OR uut_a_4_1 /= "000000000000010100011000111" OR uut_a_4_2 /= "111111111001010011110100111" OR uut_a_4_3 /= "000000000000000001000011100" OR uut_a_4_4 /= "000000000000000100001110010" OR uut_a_4_5 /= "111111111110100111010100000" OR uut_a_5_0 /= "111111111110010100111101001" OR uut_a_5_1 /= "111111111001010011110100111" OR uut_a_5_2 /= "000010001100011111100111101" OR uut_a_5_3 /= "111111111111101001110101000" OR uut_a_5_4 /= "111111111110100111010100000" OR uut_a_5_5 /= "000000011101000110011010000" THEN
              FAIL <= '1';
              FAIL_NUM <= "10101111";
              state <= "11111101";
            ELSE
              state <= "10111101";
            END IF;
            uut_rst <= '0';
          WHEN "10111101" =>
            uut_coord_shift <= "1000";
            uut_x <= "111011101010";
            uut_y <= "111101111100";
            uut_fx <= "0110010000";
            uut_fy <= "0101101101";
            uut_ft <= "1110011100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000001001011000010" OR uut_a_0_1 /= "000000010000100011110100010" OR uut_a_0_2 /= "000000000101110010011101111" OR uut_a_0_3 /= "111111111110111101011001000" OR uut_a_0_4 /= "111110001010011001001001000" OR uut_a_0_5 /= "111111010110111000111011100" OR uut_a_1_0 /= "000000000000001000010001111" OR uut_a_1_1 /= "000000001110100111100111101" OR uut_a_1_2 /= "000000000101000111000011010" OR uut_a_1_3 /= "111111111111000101001100100" OR uut_a_1_4 /= "111110011000001011001100011" OR uut_a_1_5 /= "111111011011101101010000100" OR uut_a_2_0 /= "000000000000000010111001001" OR uut_a_2_1 /= "000000000101000111000011010" OR uut_a_2_2 /= "000000000001110010010100101" OR uut_a_2_3 /= "111111111111101011011100011" OR uut_a_2_4 /= "111111011011101101010000100" OR uut_a_2_5 /= "111111110011010100000100010" OR uut_a_3_0 /= "111111111110111101011001000" OR uut_a_3_1 /= "111110001010011001001001000" OR uut_a_3_2 /= "111111010110111000111011100" OR uut_a_3_3 /= "000000000111011001000100000" OR uut_a_3_4 /= "001101000011010000000100000" OR uut_a_3_5 /= "000100100011111101111110000" OR uut_a_4_0 /= "111111111111000101001100100" OR uut_a_4_1 /= "111110011000001011001100011" OR uut_a_4_2 /= "111111011011101101010000100" OR uut_a_4_3 /= "000000000110100001101000000" OR uut_a_4_4 /= "001011100001010111101011100" OR uut_a_4_5 /= "000100000001110000001101001" OR uut_a_5_0 /= "111111111111101011011100011" OR uut_a_5_1 /= "111111011011101101010000100" OR uut_a_5_2 /= "111111110011010100000100010" OR uut_a_5_3 /= "000000000010010001111110111" OR uut_a_5_4 /= "000100000001110000001101001" OR uut_a_5_5 /= "000001011010000110010111111" THEN
              FAIL <= '1';
              FAIL_NUM <= "10110000";
              state <= "11111101";
            ELSE
              state <= "10111110";
            END IF;
            uut_rst <= '0';
          WHEN "10111110" =>
            uut_coord_shift <= "1000";
            uut_x <= "111101000110";
            uut_y <= "000001101111";
            uut_fx <= "0110100100";
            uut_fy <= "0110100011";
            uut_ft <= "0001011110";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001001000010000000" OR uut_a_0_1 /= "000000001111001111011000000" OR uut_a_0_2 /= "000000110011111011100000000" OR uut_a_0_3 /= "000000000010001101110110000" OR uut_a_0_4 /= "000000011101111010111001000" OR uut_a_0_5 /= "000001100101111100110100000" OR uut_a_1_0 /= "000000000000000111100111101" OR uut_a_1_1 /= "000000000001100110110111110" OR uut_a_1_2 /= "000000000101011110100001101" OR uut_a_1_3 /= "000000000000001110111101011" OR uut_a_1_4 /= "000000000011001001111101100" OR uut_a_1_5 /= "000000001010110000001010011" OR uut_a_2_0 /= "000000000000011001111101110" OR uut_a_2_1 /= "000000000101011110100001101" OR uut_a_2_2 /= "000000010010101010011000100" OR uut_a_2_3 /= "000000000000110010111110011" OR uut_a_2_4 /= "000000001010110000001010011" OR uut_a_2_5 /= "000000100100101000110110101" OR uut_a_3_0 /= "000000000010001101110110000" OR uut_a_3_1 /= "000000011101111010111001000" OR uut_a_3_2 /= "000001100101111100110100000" OR uut_a_3_3 /= "000000000100010110011110010" OR uut_a_3_4 /= "000000111010101111011000011" OR uut_a_3_5 /= "000011001000001001101111100" OR uut_a_4_0 /= "000000000000001110111101011" OR uut_a_4_1 /= "000000000011001001111101100" OR uut_a_4_2 /= "000000001010110000001010011" OR uut_a_4_3 /= "000000000000011101010111101" OR uut_a_4_4 /= "000000000110001100011111110" OR uut_a_4_5 /= "000000010101000111000001110" OR uut_a_5_0 /= "000000000000110010111110011" OR uut_a_5_1 /= "000000001010110000001010011" OR uut_a_5_2 /= "000000100100101000110110101" OR uut_a_5_3 /= "000000000001100100000100110" OR uut_a_5_4 /= "000000010101000111000001110" OR uut_a_5_5 /= "000001000111111011100000000" THEN
              FAIL <= '1';
              FAIL_NUM <= "10110001";
              state <= "11111101";
            ELSE
              state <= "10111111";
            END IF;
            uut_rst <= '0';
          WHEN "10111111" =>
            uut_coord_shift <= "1000";
            uut_x <= "111101010101";
            uut_y <= "000101101001";
            uut_fx <= "1111000101";
            uut_fy <= "0110011110";
            uut_ft <= "1000100010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000001001100111101010010" OR uut_a_0_1 /= "001110000011011100001110011" OR uut_a_0_2 /= "111100011101111011111111001" OR uut_a_0_3 /= "000000000001011001111100100" OR uut_a_0_4 /= "000010000011011001111000110" OR uut_a_0_5 /= "111111011110111110010010010" OR uut_a_1_0 /= "000000000111000001101110000" OR uut_a_1_1 /= "001010010001000000110111100" OR uut_a_1_2 /= "111101011010110111100100010" OR uut_a_1_3 /= "000000000001000001101100111" OR uut_a_1_4 /= "000001011111111111001010001" OR uut_a_1_5 /= "111111100111110111111111110" OR uut_a_2_0 /= "111111111110001110111101111" OR uut_a_2_1 /= "111101011010110111100100010" OR uut_a_2_2 /= "000000101001100000001111001" OR uut_a_2_3 /= "111111111111101111011111001" OR uut_a_2_4 /= "111111100111110111111111110" OR uut_a_2_5 /= "000000000110000100000100001" OR uut_a_3_0 /= "000000000001011001111100100" OR uut_a_3_1 /= "000010000011011001111000110" OR uut_a_3_2 /= "111111011110111110010010010" OR uut_a_3_3 /= "000000000000001101001001000" OR uut_a_3_4 /= "000000010011001100101001100" OR uut_a_3_5 /= "111111111011001011001100100" OR uut_a_4_0 /= "000000000001000001101100111" OR uut_a_4_1 /= "000001011111111111001010001" OR uut_a_4_2 /= "111111100111110111111111110" OR uut_a_4_3 /= "000000000000001001100110010" OR uut_a_4_4 /= "000000001110000001011111010" OR uut_a_4_5 /= "111111111100011110011011011" OR uut_a_5_0 /= "111111111111101111011111001" OR uut_a_5_1 /= "111111100111110111111111110" OR uut_a_5_2 /= "000000000110000100000100001" OR uut_a_5_3 /= "111111111111111101100101100" OR uut_a_5_4 /= "111111111100011110011011011" OR uut_a_5_5 /= "000000000000111000101100011" THEN
              FAIL <= '1';
              FAIL_NUM <= "10110010";
              state <= "11111101";
            ELSE
              state <= "11000000";
            END IF;
            uut_rst <= '0';
          WHEN "11000000" =>
            uut_coord_shift <= "1000";
            uut_x <= "000000100001";
            uut_y <= "000011011101";
            uut_fx <= "1010111000";
            uut_fy <= "1101011001";
            uut_ft <= "1011000000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000100110010010010" OR uut_a_0_1 /= "111111110001000010110111110" OR uut_a_0_2 /= "000000110010110110001111010" OR uut_a_0_3 /= "000000000000101011010100000" OR uut_a_0_4 /= "111111101111000101001100000" OR uut_a_0_5 /= "000000111001100001100100000" OR uut_a_1_0 /= "111111111111111000100001011" OR uut_a_1_1 /= "000000000010111010111100000" OR uut_a_1_2 /= "111111110110000100011010000" OR uut_a_1_3 /= "111111111111110111100010100" OR uut_a_1_4 /= "000000000011010011011111001" OR uut_a_1_5 /= "111111110100110000111100011" OR uut_a_2_0 /= "000000000000011001011011000" OR uut_a_2_1 /= "111111110110000100011010000" OR uut_a_2_2 /= "000000100001110001000001001" OR uut_a_2_3 /= "000000000000011100110000110" OR uut_a_2_4 /= "111111110100110000111100011" OR uut_a_2_5 /= "000000100110001100110010011" OR uut_a_3_0 /= "000000000000101011010100000" OR uut_a_3_1 /= "111111101111000101001100000" OR uut_a_3_2 /= "000000111001100001100100000" OR uut_a_3_3 /= "000000000000110001000000000" OR uut_a_3_4 /= "111111101100110111000000000" OR uut_a_3_5 /= "000001000001000101000000000" OR uut_a_4_0 /= "111111111111110111100010100" OR uut_a_4_1 /= "000000000011010011011111001" OR uut_a_4_2 /= "111111110100110000111100011" OR uut_a_4_3 /= "111111111111110110011011100" OR uut_a_4_4 /= "000000000011101111010000100" OR uut_a_4_5 /= "111111110011010010100001100" OR uut_a_5_0 /= "000000000000011100110000110" OR uut_a_5_1 /= "111111110100110000111100011" OR uut_a_5_2 /= "000000100110001100110010011" OR uut_a_5_3 /= "000000000000100000100010100" OR uut_a_5_4 /= "111111110011010010100001100" OR uut_a_5_5 /= "000000101011001101110100100" THEN
              FAIL <= '1';
              FAIL_NUM <= "10110011";
              state <= "11111101";
            ELSE
              state <= "11000001";
            END IF;
            uut_rst <= '0';
          WHEN "11000001" =>
            uut_coord_shift <= "1000";
            uut_x <= "111101001010";
            uut_y <= "111110011110";
            uut_fx <= "0000110010";
            uut_fy <= "1000110010";
            uut_ft <= "0000110110";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000101011101011110001" OR uut_a_0_1 /= "110000010011010001011001000" OR uut_a_0_2 /= "110101100011000101110101101" OR uut_a_0_3 /= "000000000000111011011111000" OR uut_a_0_4 /= "111101010100111110111000000" OR uut_a_0_5 /= "111110001110001001001010100" OR uut_a_1_0 /= "111111111100000100110100010" OR uut_a_1_1 /= "001011010010001001100000000" OR uut_a_1_2 /= "000111100000110001110011011" OR uut_a_1_3 /= "111111111111010101001111101" OR uut_a_1_4 /= "000001111010111010110011110" OR uut_a_1_5 /= "000001010001110101011010011" OR uut_a_2_0 /= "111111111101011000110001011" OR uut_a_2_1 /= "000111100000110001110011011" OR uut_a_2_2 /= "000101000000000101010101001" OR uut_a_2_3 /= "111111111111100011100010010" OR uut_a_2_4 /= "000001010001110101011010011" OR uut_a_2_5 /= "000000110110011110110111010" OR uut_a_3_0 /= "000000000000111011011111000" OR uut_a_3_1 /= "111101010100111110111000000" OR uut_a_3_2 /= "111110001110001001001010100" OR uut_a_3_3 /= "000000000000001010001000000" OR uut_a_3_4 /= "111111100010111001000000000" OR uut_a_3_5 /= "111111101100100111101100000" OR uut_a_4_0 /= "111111111111010101001111101" OR uut_a_4_1 /= "000001111010111010110011110" OR uut_a_4_2 /= "000001010001110101011010011" OR uut_a_4_3 /= "111111111111111000101110010" OR uut_a_4_4 /= "000000010100111011000010000" OR uut_a_4_5 /= "000000001101111011011110011" OR uut_a_5_0 /= "111111111111100011100010010" OR uut_a_5_1 /= "000001010001110101011010011" OR uut_a_5_2 /= "000000110110011110110111010" OR uut_a_5_3 /= "111111111111111011001001111" OR uut_a_5_4 /= "000000001101111011011110011" OR uut_a_5_5 /= "000000001001010001100000100" THEN
              FAIL <= '1';
              FAIL_NUM <= "10110100";
              state <= "11111101";
            ELSE
              state <= "11000010";
            END IF;
            uut_rst <= '0';
          WHEN "11000010" =>
            uut_coord_shift <= "1000";
            uut_x <= "111100011010";
            uut_y <= "111011111000";
            uut_fx <= "1011111001";
            uut_fy <= "1010011110";
            uut_ft <= "0111010011";
            uut_valid_in <= '1';
            uut_done <= '1';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000100101001000100100" OR uut_a_0_1 /= "111000011111100101001110010" OR uut_a_0_2 /= "111101001111100111010101000" OR uut_a_0_3 /= "000000000000000011110011110" OR uut_a_0_4 /= "111111111001110101110011111" OR uut_a_0_5 /= "111111111101101111010001100" OR uut_a_1_0 /= "111111111110000111111001010" OR uut_a_1_1 /= "000011000010001110110100110" OR uut_a_1_2 /= "000001000111010011111110011" OR uut_a_1_3 /= "111111111111111110011101011" OR uut_a_1_4 /= "000000000010011111010111101" OR uut_a_1_5 /= "000000000000111010100000110" OR uut_a_2_0 /= "111111111111010011111001110" OR uut_a_2_1 /= "000001000111010011111110011" OR uut_a_2_2 /= "000000011010001011101010011" OR uut_a_2_3 /= "111111111111111111011011110" OR uut_a_2_4 /= "000000000000111010100000110" OR uut_a_2_5 /= "000000000000010101011110111" OR uut_a_3_0 /= "000000000000000011110011110" OR uut_a_3_1 /= "111111111001110101110011111" OR uut_a_3_2 /= "111111111101101111010001100" OR uut_a_3_3 /= "000000000000000000000011001" OR uut_a_3_4 /= "111111111111111010111100100" OR uut_a_3_5 /= "111111111111111110001001010" OR uut_a_4_0 /= "111111111111111110011101011" OR uut_a_4_1 /= "000000000010011111010111101" OR uut_a_4_2 /= "000000000000111010100000110" OR uut_a_4_3 /= "111111111111111111111110101" OR uut_a_4_4 /= "000000000000000010000010110" OR uut_a_4_5 /= "000000000000000000110000000" OR uut_a_5_0 /= "111111111111111111011011110" OR uut_a_5_1 /= "000000000000111010100000110" OR uut_a_5_2 /= "000000000000010101011110111" OR uut_a_5_3 /= "111111111111111111111111100" OR uut_a_5_4 /= "000000000000000000110000000" OR uut_a_5_5 /= "000000000000000000010001101" THEN
              FAIL <= '1';
              FAIL_NUM <= "10110101";
              state <= "11111101";
            ELSE
              state <= "11000011";
            END IF;
            uut_rst <= '0';
          WHEN "11000011" =>
            uut_coord_shift <= "1000";
            uut_x <= "000110111110";
            uut_y <= "000101000110";
            uut_fx <= "0011101010";
            uut_fy <= "1010110100";
            uut_ft <= "1101110001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000101110011010010000" OR uut_a_0_1 /= "110100001000000010001010000" OR uut_a_0_2 /= "001101001100000101011011000" OR uut_a_0_3 /= "000000000001011100110100100" OR uut_a_0_4 /= "111101000010000000100010100" OR uut_a_0_5 /= "000011010011000001010110110" OR uut_a_1_0 /= "111111111101000010000000100" OR uut_a_1_1 /= "000110000100111000111001011" OR uut_a_1_2 /= "111001010000000100001110011" OR uut_a_1_3 /= "111111111111010000100000001" OR uut_a_1_4 /= "000001100001001110001110010" OR uut_a_1_5 /= "111110010100000001000011100" OR uut_a_2_0 /= "000000000011010011000001010" OR uut_a_2_1 /= "111001010000000100001110011" OR uut_a_2_2 /= "000111011111101111100101001" OR uut_a_2_3 /= "000000000000110100110000010" OR uut_a_2_4 /= "111110010100000001000011100" OR uut_a_2_5 /= "000001110111111011111001010" OR uut_a_3_0 /= "000000000001011100110100100" OR uut_a_3_1 /= "111101000010000000100010100" OR uut_a_3_2 /= "000011010011000001010110110" OR uut_a_3_3 /= "000000000000010111001101001" OR uut_a_3_4 /= "111111010000100000001000101" OR uut_a_3_5 /= "000000110100110000010101101" OR uut_a_4_0 /= "111111111111010000100000001" OR uut_a_4_1 /= "000001100001001110001110010" OR uut_a_4_2 /= "111110010100000001000011100" OR uut_a_4_3 /= "111111111111110100001000000" OR uut_a_4_4 /= "000000011000010011100011100" OR uut_a_4_5 /= "111111100101000000010000111" OR uut_a_5_0 /= "000000000000110100110000010" OR uut_a_5_1 /= "111110010100000001000011100" OR uut_a_5_2 /= "000001110111111011111001010" OR uut_a_5_3 /= "000000000000001101001100000" OR uut_a_5_4 /= "111111100101000000010000111" OR uut_a_5_5 /= "000000011101111110111110010" THEN
              FAIL <= '1';
              FAIL_NUM <= "10110110";
              state <= "11111101";
            ELSE
              state <= "11000100";
            END IF;
            uut_rst <= '0';
          WHEN "11000100" =>
            uut_coord_shift <= "1000";
            uut_x <= "111011000010";
            uut_y <= "111000000010";
            uut_fx <= "1101000100";
            uut_fy <= "0011001100";
            uut_ft <= "0010000000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000011000101100000100" OR uut_a_0_1 /= "111001000110101100011000100" OR uut_a_0_2 /= "110011101101000011100000100" OR uut_a_0_3 /= "000000000011100011010100100" OR uut_a_0_4 /= "111000000100000101001100100" OR uut_a_0_5 /= "110001110110010001010100100" OR uut_a_1_0 /= "111111111110010001101011000" OR uut_a_1_1 /= "000011110110100000101101010" OR uut_a_1_2 /= "000110110111100101010010100" OR uut_a_1_3 /= "111111111110000001000001010" OR uut_a_1_4 /= "000100011011101110000110010" OR uut_a_1_5 /= "000111111001111011110100110" OR uut_a_2_0 /= "111111111100111011010000111" OR uut_a_2_1 /= "000110110111100101010010100" OR uut_a_2_2 /= "001100001111110111110000011" OR uut_a_2_3 /= "111111111100011101100100010" OR uut_a_2_4 /= "000111111001111011110100110" OR uut_a_2_5 /= "001110000110001100001111110" OR uut_a_3_0 /= "000000000011100011010100100" OR uut_a_3_1 /= "111000000100000101001100100" OR uut_a_3_2 /= "110001110110010001010100100" OR uut_a_3_3 /= "000000000100000101101000100" OR uut_a_3_4 /= "110110110111011010100000100" OR uut_a_3_5 /= "101111101101100011101000100" OR uut_a_4_0 /= "111111111110000001000001010" OR uut_a_4_1 /= "000100011011101110000110010" OR uut_a_4_2 /= "000111111001111011110100110" OR uut_a_4_3 /= "111111111101101101110110101" OR uut_a_4_4 /= "000101000110100010111100010" OR uut_a_4_5 /= "001001000110010011010110001" OR uut_a_5_0 /= "111111111100011101100100010" OR uut_a_5_1 /= "000111111001111011110100110" OR uut_a_5_2 /= "001110000110001100001111110" OR uut_a_5_3 /= "111111111011111011011000111" OR uut_a_5_4 /= "001001000110010011010110001" OR uut_a_5_5 /= "010000001110010111110000011" THEN
              FAIL <= '1';
              FAIL_NUM <= "10110111";
              state <= "11111101";
            ELSE
              state <= "11000101";
            END IF;
            uut_rst <= '0';
          WHEN "11000101" =>
            uut_coord_shift <= "1000";
            uut_x <= "000000101100";
            uut_y <= "111111000010";
            uut_fx <= "1100100110";
            uut_fy <= "0000000010";
            uut_ft <= "0100001100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000010011111011001" OR uut_a_0_1 /= "111111001100010100101001010" OR uut_a_0_2 /= "111111000110011010000101111" OR uut_a_0_3 /= "000000000001010001000100111" OR uut_a_0_4 /= "111100101101101101010110110" OR uut_a_0_5 /= "111100010101101000111010001" OR uut_a_1_0 /= "111111111111110011000101001" OR uut_a_1_1 /= "000000100001100000100111010" OR uut_a_1_2 /= "000000100101010110000101001" OR uut_a_1_3 /= "111111111111001011011011010" OR uut_a_1_4 /= "000010001000010111000101101" OR uut_a_1_5 /= "000010010111111101111110010" OR uut_a_2_0 /= "111111111111110001100110100" OR uut_a_2_1 /= "000000100101010110000101001" OR uut_a_2_2 /= "000000101001100111101001010" OR uut_a_2_3 /= "111111111111000101011010001" OR uut_a_2_4 /= "000010010111111101111110010" OR uut_a_2_5 /= "000010101001010111001011111" OR uut_a_3_0 /= "000000000001010001000100111" OR uut_a_3_1 /= "111100101101101101010110110" OR uut_a_3_2 /= "111100010101101000111010001" OR uut_a_3_3 /= "000000000101001001111011001" OR uut_a_3_4 /= "110010101000010000101001010" OR uut_a_3_5 /= "110001000110010100000101111" OR uut_a_4_0 /= "111111111111001011011011010" OR uut_a_4_1 /= "000010001000010111000101101" OR uut_a_4_2 /= "000010010111111101111110010" OR uut_a_4_3 /= "111111111100101010000100001" OR uut_a_4_4 /= "001000101010111001001101010" OR uut_a_4_5 /= "001001101010011001111110001" OR uut_a_5_0 /= "111111111111000101011010001" OR uut_a_5_1 /= "000010010111111101111110010" OR uut_a_5_2 /= "000010101001010111001011111" OR uut_a_5_3 /= "111111111100010001100101000" OR uut_a_5_4 /= "001001101010011001111110001" OR uut_a_5_5 /= "001010110001001011111110110" THEN
              FAIL <= '1';
              FAIL_NUM <= "10111000";
              state <= "11111101";
            ELSE
              state <= "11000110";
            END IF;
            uut_rst <= '0';
          WHEN "11000110" =>
            uut_coord_shift <= "1000";
            uut_x <= "000100001100";
            uut_y <= "000001001101";
            uut_fx <= "0011111110";
            uut_fy <= "0010010101";
            uut_ft <= "1001111110";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000011111100000001" OR uut_a_0_1 /= "111110111001110110111110001" OR uut_a_0_2 /= "111111111011110100001110111" OR uut_a_0_3 /= "111111111111111010000011000" OR uut_a_0_4 /= "000000001101010000010100100" OR uut_a_0_5 /= "000000000000110010100110100" OR uut_a_1_0 /= "111111111111101110011101101" OR uut_a_1_1 /= "000000100111000010110001101" OR uut_a_1_2 /= "000000000010010101000011001" OR uut_a_1_3 /= "000000000000000011010100000" OR uut_a_1_4 /= "111111111000100111110010100" OR uut_a_1_5 /= "111111111111100011110101010" OR uut_a_2_0 /= "111111111111111110111101000" OR uut_a_2_1 /= "000000000010010101000011001" OR uut_a_2_2 /= "000000000000001000111001000" OR uut_a_2_3 /= "000000000000000000001100101" OR uut_a_2_4 /= "111111111111100011110101010" OR uut_a_2_5 /= "111111111111111110010100011" OR uut_a_3_0 /= "111111111111111010000011000" OR uut_a_3_1 /= "000000001101010000010100100" OR uut_a_3_2 /= "000000000000110010100110100" OR uut_a_3_3 /= "000000000000000001001000000" OR uut_a_3_4 /= "111111111101011111101100000" OR uut_a_3_5 /= "111111111111110110011100000" OR uut_a_4_0 /= "000000000000000011010100000" OR uut_a_4_1 /= "111111111000100111110010100" OR uut_a_4_2 /= "111111111111100011110101010" OR uut_a_4_3 /= "111111111111111111010111111" OR uut_a_4_4 /= "000000000001011001001111001" OR uut_a_4_5 /= "000000000000000101010100101" OR uut_a_5_0 /= "000000000000000000001100101" OR uut_a_5_1 /= "111111111111100011110101010" OR uut_a_5_2 /= "111111111111111110010100011" OR uut_a_5_3 /= "111111111111111111111101100" OR uut_a_5_4 /= "000000000000000101010100101" OR uut_a_5_5 /= "000000000000000000010100010" THEN
              FAIL <= '1';
              FAIL_NUM <= "10111001";
              state <= "11111101";
            ELSE
              state <= "11000111";
            END IF;
            uut_rst <= '0';
          WHEN "11000111" =>
            uut_coord_shift <= "1000";
            uut_x <= "000000000100";
            uut_y <= "111101100100";
            uut_fx <= "1001011110";
            uut_fy <= "1010010111";
            uut_ft <= "1011001011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000011011001111000100" OR uut_a_0_1 /= "110100001111100111111001100" OR uut_a_0_2 /= "111110010001010110110011110" OR uut_a_0_3 /= "000000000100111100011000110" OR uut_a_0_4 /= "101110111011011110100010010" OR uut_a_0_5 /= "111101011111010101011011101" OR uut_a_1_0 /= "111111111101000011111001111" OR uut_a_1_1 /= "001010001001100000110011100" OR uut_a_1_2 /= "000001011111100001000011110" OR uut_a_1_3 /= "111111111011101110110111101" OR uut_a_1_4 /= "001110101111001001111000111" OR uut_a_1_5 /= "000010001010101100101111111" OR uut_a_2_0 /= "111111111111100100010101101" OR uut_a_2_1 /= "000001011111100001000011110" OR uut_a_2_2 /= "000000001110000010111110101" OR uut_a_2_3 /= "111111111111010111110101010" OR uut_a_2_4 /= "000010001010101100101111111" OR uut_a_2_5 /= "000000010100011001011001110" OR uut_a_3_0 /= "000000000100111100011000110" OR uut_a_3_1 /= "101110111011011110100010010" OR uut_a_3_2 /= "111101011111010101011011101" OR uut_a_3_3 /= "000000000111001011011011001" OR uut_a_3_4 /= "100111001101100011010101011" OR uut_a_3_5 /= "111100010110101100101110011" OR uut_a_4_0 /= "111111111011101110110111101" OR uut_a_4_1 /= "001110101111001001111000111" OR uut_a_4_2 /= "000010001010101100101111111" OR uut_a_4_3 /= "111111111001110011011000110" OR uut_a_4_4 /= "010101011001100011001111110" OR uut_a_4_5 /= "000011001001011001111000111" OR uut_a_5_0 /= "111111111111010111110101010" OR uut_a_5_1 /= "000010001010101100101111111" OR uut_a_5_2 /= "000000010100011001011001110" OR uut_a_5_3 /= "111111111111000101101011001" OR uut_a_5_4 /= "000011001001011001111000111" OR uut_a_5_5 /= "000000011101100111100100100" THEN
              FAIL <= '1';
              FAIL_NUM <= "10111010";
              state <= "11111101";
            ELSE
              state <= "11001000";
            END IF;
            uut_rst <= '0';
          WHEN "11001000" =>
            uut_coord_shift <= "1001";
            uut_x <= "000101100000";
            uut_y <= "111101110100";
            uut_fx <= "0011000111";
            uut_fy <= "1100000111";
            uut_ft <= "1000001010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000010001101010101001" OR uut_a_0_1 /= "111110110001100110110010000" OR uut_a_0_2 /= "001000001001001001111001100" OR uut_a_0_3 /= "111111111011110111001101000" OR uut_a_0_4 /= "000010010010111000010010100" OR uut_a_0_5 /= "110000101111100011111100000" OR uut_a_1_0 /= "111111111111101100011001101" OR uut_a_1_1 /= "000000001010110111101111110" OR uut_a_1_2 /= "111110110111101110110000001" OR uut_a_1_3 /= "000000000000100100101110000" OR uut_a_1_4 /= "111111101011101000011100011" OR uut_a_1_5 /= "000010000111011001111001000" OR uut_a_2_0 /= "000000000010000010010010011" OR uut_a_2_1 /= "111110110111101110110000001" OR uut_a_2_2 /= "000111100000011100001000000" OR uut_a_2_3 /= "111111111100001011111000111" OR uut_a_2_4 /= "000010000111011001111001000" OR uut_a_2_5 /= "110001111011110110001000010" OR uut_a_3_0 /= "111111111011110111001101000" OR uut_a_3_1 /= "000010010010111000010010100" OR uut_a_3_2 /= "110000101111100011111100000" OR uut_a_3_3 /= "000000000111110000001000000" OR uut_a_3_4 /= "111011101100110011100100000" OR uut_a_3_5 /= "011100100101011101100000000" OR uut_a_4_0 /= "000000000000100100101110000" OR uut_a_4_1 /= "111111101011101000011100011" OR uut_a_4_2 /= "000010000111011001111001000" OR uut_a_4_3 /= "111111111110111011001100111" OR uut_a_4_4 /= "000000100110001010010110011" OR uut_a_4_5 /= "111100000010010011100010001" OR uut_a_5_0 /= "111111111100001011111000111" OR uut_a_5_1 /= "000010000111011001111001000" OR uut_a_5_2 /= "110001111011110110001000010" OR uut_a_5_3 /= "000000000111001001010111011" OR uut_a_5_4 /= "111100000010010011100010001" OR uut_a_5_5 /= "011010010110100010001100100" THEN
              FAIL <= '1';
              FAIL_NUM <= "10111011";
              state <= "11111101";
            ELSE
              state <= "11001001";
            END IF;
            uut_rst <= '0';
          WHEN "11001001" =>
            uut_coord_shift <= "1001";
            uut_x <= "000001000010";
            uut_y <= "111000111101";
            uut_fx <= "0111001001";
            uut_fy <= "0110100000";
            uut_ft <= "1110010010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000101101100100" OR uut_a_0_1 /= "000000001001010110000000100" OR uut_a_0_2 /= "000000000110100101011101000" OR uut_a_0_3 /= "111111111111100001100001010" OR uut_a_0_4 /= "111111001101111111100011010" OR uut_a_0_5 /= "111111011100110000011100100" OR uut_a_1_0 /= "000000000000000010010101100" OR uut_a_1_1 /= "000000000011110101010001101" OR uut_a_1_2 /= "000000000010101100110111001" OR uut_a_1_3 /= "111111111111110011011111111" OR uut_a_1_4 /= "111111101011011111010100001" OR uut_a_1_5 /= "111111110001100010110111101" OR uut_a_2_0 /= "000000000000000001101001010" OR uut_a_2_1 /= "000000000010101100110111001" OR uut_a_2_2 /= "000000000001111001110100111" OR uut_a_2_3 /= "111111111111110111001100000" OR uut_a_2_4 /= "111111110001100010110111101" OR uut_a_2_5 /= "111111110101110100000000001" OR uut_a_3_0 /= "111111111111100001100001010" OR uut_a_3_1 /= "111111001101111111100011010" OR uut_a_3_2 /= "111111011100110000011100100" OR uut_a_3_3 /= "000000000010100011001000001" OR uut_a_3_4 /= "000100001011101000010101001" OR uut_a_3_5 /= "000010111100100111011001010" OR uut_a_4_0 /= "111111111111110011011111111" OR uut_a_4_1 /= "111111101011011111010100001" OR uut_a_4_2 /= "111111110001100010110111101" OR uut_a_4_3 /= "000000000001000010111010000" OR uut_a_4_4 /= "000001101101110001010010101" OR uut_a_4_5 /= "000001001101010111001010000" OR uut_a_5_0 /= "111111111111110111001100000" OR uut_a_5_1 /= "111111110001100010110111101" OR uut_a_5_2 /= "111111110101110100000000001" OR uut_a_5_3 /= "000000000000101111001001110" OR uut_a_5_4 /= "000001001101010111001010000" OR uut_a_5_5 /= "000000110110100001011000110" THEN
              FAIL <= '1';
              FAIL_NUM <= "10111100";
              state <= "11111101";
            ELSE
              state <= "11001010";
            END IF;
            uut_rst <= '0';
          WHEN "11001010" =>
            uut_coord_shift <= "1001";
            uut_x <= "110000110011";
            uut_y <= "000101011111";
            uut_fx <= "0101011001";
            uut_fy <= "0111100011";
            uut_ft <= "1000111010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000100111000100000000" OR uut_a_0_1 /= "110101011001010010100000000" OR uut_a_0_2 /= "111010111101101111000000000" OR uut_a_0_3 /= "000000000100011101001010000" OR uut_a_0_4 /= "110110010100101011010010000" OR uut_a_0_5 /= "111011011001111011101100000" OR uut_a_1_0 /= "111111111101010110010100101" OR uut_a_1_1 /= "000101110000100001001101001" OR uut_a_1_2 /= "000010101110111110101110110" OR uut_a_1_3 /= "111111111101100101001010110" OR uut_a_1_4 /= "000101010000010001011111111" OR uut_a_1_5 /= "000010011111101010110101110" OR uut_a_2_0 /= "111111111110101111011011110" OR uut_a_2_1 /= "000010101110111110101110110" OR uut_a_2_2 /= "000001010011000101011000100" OR uut_a_2_3 /= "111111111110110110011110111" OR uut_a_2_4 /= "000010011111101010110101110" OR uut_a_2_5 /= "000001001011110100000111001" OR uut_a_3_0 /= "000000000100011101001010000" OR uut_a_3_1 /= "110110010100101011010010000" OR uut_a_3_2 /= "111011011001111011101100000" OR uut_a_3_3 /= "000000000100000100001101001" OR uut_a_3_4 /= "110111001010110111011111101" OR uut_a_3_5 /= "111011110011101010011101110" OR uut_a_4_0 /= "111111111101100101001010110" OR uut_a_4_1 /= "000101010000010001011111111" OR uut_a_4_2 /= "000010011111101010110101110" OR uut_a_4_3 /= "111111111101110010101101110" OR uut_a_4_4 /= "000100110010110110010111100" OR uut_a_4_5 /= "000010010001101100101100010" OR uut_a_5_0 /= "111111111110110110011110111" OR uut_a_5_1 /= "000010011111101010110101110" OR uut_a_5_2 /= "000001001011110100000111001" OR uut_a_5_3 /= "111111111110111100111010100" OR uut_a_5_4 /= "000010010001101100101100010" OR uut_a_5_5 /= "000001000101001011100011010" THEN
              FAIL <= '1';
              FAIL_NUM <= "10111101";
              state <= "11111101";
            ELSE
              state <= "11001011";
            END IF;
            uut_rst <= '0';
          WHEN "11001011" =>
            uut_coord_shift <= "1001";
            uut_x <= "111110011011";
            uut_y <= "000010101000";
            uut_fx <= "0010111111";
            uut_fy <= "0011100001";
            uut_ft <= "0010011010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000101011000100010000" OR uut_a_0_1 /= "111000001011010110100110000" OR uut_a_0_2 /= "000100101010110001011111000" OR uut_a_0_3 /= "000000000101010111101101100" OR uut_a_0_4 /= "111000001100100010111000100" OR uut_a_0_5 /= "000100101010000011111101010" OR uut_a_1_0 /= "111111111110000010110101101" OR uut_a_1_1 /= "000010110101111000000010101" OR uut_a_1_2 /= "111110010011011101100001011" OR uut_a_1_3 /= "111111111110000011001000101" OR uut_a_1_4 /= "000010110101011100010100111" OR uut_a_1_5 /= "111110010011101110000011111" OR uut_a_2_0 /= "000000000001001010101100010" OR uut_a_2_1 /= "111110010011011101100001011" OR uut_a_2_2 /= "000001000000110001011110100" OR uut_a_2_3 /= "000000000001001010100000111" OR uut_a_2_4 /= "111110010011101110000011111" OR uut_a_2_5 /= "000001000000100111100110111" OR uut_a_3_0 /= "000000000101010111101101100" OR uut_a_3_1 /= "111000001100100010111000100" OR uut_a_3_2 /= "000100101010000011111101010" OR uut_a_3_3 /= "000000000101010110111001001" OR uut_a_3_4 /= "111000001101101110111111011" OR uut_a_3_5 /= "000100101001010110100010011" OR uut_a_4_0 /= "111111111110000011001000101" OR uut_a_4_1 /= "000010110101011100010100111" OR uut_a_4_2 /= "111110010011101110000011111" OR uut_a_4_3 /= "111111111110000011011011101" OR uut_a_4_4 /= "000010110101000000101011011" OR uut_a_4_5 /= "111110010011111110100011111" OR uut_a_5_0 /= "000000000001001010100000111" OR uut_a_5_1 /= "111110010011101110000011111" OR uut_a_5_2 /= "000001000000100111100110111" OR uut_a_5_3 /= "000000000001001010010101101" OR uut_a_5_4 /= "111110010011111110100011111" OR uut_a_5_5 /= "000001000000011101110000101" THEN
              FAIL <= '1';
              FAIL_NUM <= "10111110";
              state <= "11111101";
            ELSE
              state <= "11001100";
            END IF;
            uut_rst <= '0';
          WHEN "11001100" =>
            uut_coord_shift <= "1001";
            uut_x <= "000111010000";
            uut_y <= "111011111110";
            uut_fx <= "0001010100";
            uut_fy <= "1001110111";
            uut_ft <= "1000111011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000110110011001" OR uut_a_0_1 /= "111111110110111010101100110" OR uut_a_0_2 /= "000000010011001011001100000" OR uut_a_0_3 /= "111111111111010000010010110" OR uut_a_0_4 /= "000000111111101110111100111" OR uut_a_0_5 /= "111101111001011100111000011" OR uut_a_1_0 /= "111111111111111101101110101" OR uut_a_1_1 /= "000000000011000010001001010" OR uut_a_1_2 /= "111111111001100110001000110" OR uut_a_1_3 /= "000000000000001111111011101" OR uut_a_1_4 /= "111111101010101101101100011" OR uut_a_1_5 /= "000000101100111011111110101" OR uut_a_2_0 /= "000000000000000100110010110" OR uut_a_2_1 /= "111111111001100110001000110" OR uut_a_2_2 /= "000000001101100001010000111" OR uut_a_2_3 /= "111111111111011110010111001" OR uut_a_2_4 /= "000000101100111011111110101" OR uut_a_2_5 /= "111110100001001000011111001" OR uut_a_3_0 /= "111111111111010000010010110" OR uut_a_3_1 /= "000000111111101110111100111" OR uut_a_3_2 /= "111101111001011100111000011" OR uut_a_3_3 /= "000000000101001110110000100" OR uut_a_3_4 /= "111001000000110010001101010" OR uut_a_3_5 /= "001110110000000111110010010" OR uut_a_4_0 /= "000000000000001111111011101" OR uut_a_4_1 /= "111111101010101101101100011" OR uut_a_4_2 /= "000000101100111011111110101" OR uut_a_4_3 /= "111111111110010000001100100" OR uut_a_4_4 /= "000010010101010111001110110" OR uut_a_4_5 /= "111011000100101011011001100" OR uut_a_5_0 /= "111111111111011110010111001" OR uut_a_5_1 /= "000000101100111011111110101" OR uut_a_5_2 /= "111110100001001000011111001" OR uut_a_5_3 /= "000000000011101100000001111" OR uut_a_5_4 /= "111011000100101011011001100" OR uut_a_5_5 /= "001010011001101011011111010" THEN
              FAIL <= '1';
              FAIL_NUM <= "10111111";
              state <= "11111101";
            ELSE
              state <= "11001101";
            END IF;
            uut_rst <= '0';
          WHEN "11001101" =>
            uut_coord_shift <= "1001";
            uut_x <= "001111010110";
            uut_y <= "111001001000";
            uut_fx <= "0001100001";
            uut_fy <= "0111011001";
            uut_ft <= "1010111110";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000011010010001000000" OR uut_a_0_1 /= "000000110110001011000100000" OR uut_a_0_2 /= "000101101010110010110100000" OR uut_a_0_3 /= "000000000001101010111111000" OR uut_a_0_4 /= "000000011011100101001111100" OR uut_a_0_5 /= "000010111000101101110001100" OR uut_a_1_0 /= "000000000000001101100010110" OR uut_a_1_1 /= "000000000011011111011101101" OR uut_a_1_2 /= "000000010111011000100001100" OR uut_a_1_3 /= "000000000000000110111001010" OR uut_a_1_4 /= "000000000001110001110001100" OR uut_a_1_5 /= "000000001011111001111100110" OR uut_a_2_0 /= "000000000001011010101100101" OR uut_a_2_1 /= "000000010111011000100001100" OR uut_a_2_2 /= "000010011100100110001011101" OR uut_a_2_3 /= "000000000000101110001011011" OR uut_a_2_4 /= "000000001011111001111100110" OR uut_a_2_5 /= "000001001111101110110000011" OR uut_a_3_0 /= "000000000001101010111111000" OR uut_a_3_1 /= "000000011011100101001111100" OR uut_a_3_2 /= "000010111000101101110001100" OR uut_a_3_3 /= "000000000000110110011110001" OR uut_a_3_4 /= "000000001110000010110001000" OR uut_a_3_5 /= "000001011110000011000000110" OR uut_a_4_0 /= "000000000000000110111001010" OR uut_a_4_1 /= "000000000001110001110001100" OR uut_a_4_2 /= "000000001011111001111100110" OR uut_a_4_3 /= "000000000000000011100000101" OR uut_a_4_4 /= "000000000000111001111011011" OR uut_a_4_5 /= "000000000110000011111100011" OR uut_a_5_0 /= "000000000000101110001011011" OR uut_a_5_1 /= "000000001011111001111100110" OR uut_a_5_2 /= "000001001111101110110000011" OR uut_a_5_3 /= "000000000000010111100000110" OR uut_a_5_4 /= "000000000110000011111100011" OR uut_a_5_5 /= "000000101000100110000011001" THEN
              FAIL <= '1';
              FAIL_NUM <= "11000000";
              state <= "11111101";
            ELSE
              state <= "11001110";
            END IF;
            uut_rst <= '0';
          WHEN "11001110" =>
            uut_coord_shift <= "1001";
            uut_x <= "110110001100";
            uut_y <= "111010111100";
            uut_fx <= "0110111011";
            uut_fy <= "1110010000";
            uut_ft <= "1100011000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000100111000100" OR uut_a_0_1 /= "111111111001000011101010100" OR uut_a_0_2 /= "111111111100010000101111100" OR uut_a_0_3 /= "111111111111010010111000100" OR uut_a_0_4 /= "000001000000001001101010100" OR uut_a_0_5 /= "000000100010100010101111100" OR uut_a_1_0 /= "111111111111111110010000111" OR uut_a_1_1 /= "000000000010011101111100101" OR uut_a_1_2 /= "000000000001010101000011000" OR uut_a_1_3 /= "000000000000010000000010011" OR uut_a_1_4 /= "111111101001001100100100001" OR uut_a_1_5 /= "111111110011101110001001100" OR uut_a_2_0 /= "111111111111111111000100001" OR uut_a_2_1 /= "000000000001010101000011000" OR uut_a_2_2 /= "000000000000101101110010111" OR uut_a_2_3 /= "000000000000001000101000101" OR uut_a_2_4 /= "111111110011101110001001100" OR uut_a_2_5 /= "111111111001011000110110011" OR uut_a_3_0 /= "111111111111010010111000100" OR uut_a_3_1 /= "000001000000001001101010100" OR uut_a_3_2 /= "000000100010100010101111100" OR uut_a_3_3 /= "000000000110100000111000100" OR uut_a_3_4 /= "110110101111001111101010100" OR uut_a_3_5 /= "111011000000110100101111100" OR uut_a_4_0 /= "000000000000010000000010011" OR uut_a_4_1 /= "111111101001001100100100001" OR uut_a_4_2 /= "111111110011101110001001100" OR uut_a_4_3 /= "111111111101101011110011111" OR uut_a_4_4 /= "000011010010101101001011101" OR uut_a_4_5 /= "000001110001011101010000000" OR uut_a_5_0 /= "000000000000001000101000101" OR uut_a_5_1 /= "111111110011101110001001100" OR uut_a_5_2 /= "111111111001011000110110011" OR uut_a_5_3 /= "111111111110110000001101001" OR uut_a_5_4 /= "000001110001011101010000000" OR uut_a_5_5 /= "000000111101000101111001111" THEN
              FAIL <= '1';
              FAIL_NUM <= "11000001";
              state <= "11111101";
            ELSE
              state <= "11001111";
            END IF;
            uut_rst <= '0';
          WHEN "11001111" =>
            uut_coord_shift <= "1001";
            uut_x <= "110100111000";
            uut_y <= "111100101110";
            uut_fx <= "1110000000";
            uut_fy <= "1010000110";
            uut_ft <= "1110111101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '1' OR uut_a_0_0 /= "000000000010000111000110001" OR uut_a_0_1 /= "111100001101001111111111101" OR uut_a_0_2 /= "111011101001010111010111100" OR uut_a_0_3 /= "000000000010110101110101110" OR uut_a_0_4 /= "111010111001010000011010110" OR uut_a_0_5 /= "111010001000111101001001000" OR uut_a_1_0 /= "111111111111000011010011111" OR uut_a_1_1 /= "000001101101000011000100001" OR uut_a_1_2 /= "000001111101001010110000001" OR uut_a_1_3 /= "111111111110101110010100000" OR uut_a_1_4 /= "000010010010110001110111111" OR uut_a_1_5 /= "000010101000011110100010001" OR uut_a_2_0 /= "111111111110111010010101110" OR uut_a_2_1 /= "000001111101001010110000001" OR uut_a_2_2 /= "000010001111101010111100111" OR uut_a_2_3 /= "111111111110100010001111010" OR uut_a_2_4 /= "000010101000011110100010001" OR uut_a_2_5 /= "000011000001011000011110010" OR uut_a_3_0 /= "000000000010110101110101110" OR uut_a_3_1 /= "111010111001010000011010110" OR uut_a_3_2 /= "111010001000111101001001000" OR uut_a_3_3 /= "000000000011110100110000100" OR uut_a_3_4 /= "111001001000001100110110100" OR uut_a_3_5 /= "111000000111001011111110000" OR uut_a_4_0 /= "111111111110101110010100000" OR uut_a_4_1 /= "000010010010110001110111111" OR uut_a_4_2 /= "000010101000011110100010001" OR uut_a_4_3 /= "111111111110010010000011001" OR uut_a_4_4 /= "000011000101100100001110100" OR uut_a_4_5 /= "000011100010110001010111111" OR uut_a_5_0 /= "111111111110100010001111010" OR uut_a_5_1 /= "000010101000011110100010001" OR uut_a_5_2 /= "000011000001011000011110010" OR uut_a_5_3 /= "111111111110000001110010111" OR uut_a_5_4 /= "000011100010110001010111111" OR uut_a_5_5 /= "000100000100010010110101000" THEN
              FAIL <= '1';
              FAIL_NUM <= "11000010";
              state <= "11111101";
            ELSE
              state <= "11010000";
            END IF;
            uut_rst <= '0';
          WHEN "11010000" =>
            uut_coord_shift <= "1001";
            uut_x <= "110010111100";
            uut_y <= "000011101010";
            uut_fx <= "1000001011";
            uut_fy <= "0001001011";
            uut_ft <= "0100101001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001101010111100100" OR uut_a_0_1 /= "000101110100101000110011100" OR uut_a_0_2 /= "000100010000011000000101100" OR uut_a_0_3 /= "111111111101101000010001000" OR uut_a_0_4 /= "110111101111010011001111000" OR uut_a_0_5 /= "111001111101100011010011000" OR uut_a_1_0 /= "000000000001011101001010001" OR uut_a_1_1 /= "000101000100100110100010110" OR uut_a_1_2 /= "000011101101010000111110110" OR uut_a_1_3 /= "111111111101111011110100110" OR uut_a_1_4 /= "111000110011011101000000010" OR uut_a_1_5 /= "111010101111010111011111110" OR uut_a_2_0 /= "000000000001000100000110000" OR uut_a_2_1 /= "000011101101010000111110110" OR uut_a_2_2 /= "000010101101011011010101100" OR uut_a_2_3 /= "111111111110011111011000110" OR uut_a_2_4 /= "111010101111010111011111110" OR uut_a_2_5 /= "111100001001111100001110010" OR uut_a_3_0 /= "111111111101101000010001000" OR uut_a_3_1 /= "110111101111010011001111000" OR uut_a_3_2 /= "111001111101100011010011000" OR uut_a_3_3 /= "000000000011010111010010000" OR uut_a_3_4 /= "001011101110000111101110000" OR uut_a_3_5 /= "001000100100010010110110000" OR uut_a_4_0 /= "111111111101111011110100110" OR uut_a_4_1 /= "111000110011011101000000010" OR uut_a_4_2 /= "111010101111010111011111110" OR uut_a_4_3 /= "000000000010111011100001111" OR uut_a_4_4 /= "001010001101011011001110010" OR uut_a_4_5 /= "000111011101100111011010100" OR uut_a_5_0 /= "111111111110011111011000110" OR uut_a_5_1 /= "111010101111010111011111110" OR uut_a_5_2 /= "111100001001111100001110010" OR uut_a_5_3 /= "000000000010001001000100101" OR uut_a_5_4 /= "000111011101100111011010100" OR uut_a_5_5 /= "000101011101000110111111111" THEN
              FAIL <= '1';
              FAIL_NUM <= "11000011";
              state <= "11111101";
            ELSE
              state <= "11010001";
            END IF;
            uut_rst <= '0';
          WHEN "11010001" =>
            uut_coord_shift <= "1001";
            uut_x <= "110111100011";
            uut_y <= "111110010110";
            uut_fx <= "0001000111";
            uut_fy <= "1000111111";
            uut_ft <= "1111111100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001000101000010000" OR uut_a_0_1 /= "111101010100100000000010000" OR uut_a_0_2 /= "111011101100111101000010000" OR uut_a_0_3 /= "111111111110110101000110000" OR uut_a_0_4 /= "000010111010000110000110000" OR uut_a_0_5 /= "000100101010011101000110000" OR uut_a_1_0 /= "111111111111010101001000000" OR uut_a_1_1 /= "000001101010100001000110110" OR uut_a_1_2 /= "000010101010110101000110000" OR uut_a_1_3 /= "000000000000101110100001100" OR uut_a_1_4 /= "111110001100011010101101110" OR uut_a_1_5 /= "111101000110101000011011100" OR uut_a_2_0 /= "111111111110111011001111010" OR uut_a_2_1 /= "000010101010110101000110000" OR uut_a_2_2 /= "000100010001111110001101010" OR uut_a_2_3 /= "000000000001001010100111010" OR uut_a_2_4 /= "111101000110101000011011100" OR uut_a_2_5 /= "111011010110101101100001010" OR uut_a_3_0 /= "111111111110110101000110000" OR uut_a_3_1 /= "000010111010000110000110000" OR uut_a_3_2 /= "000100101010011101000110000" OR uut_a_3_3 /= "000000000001010001010010000" OR uut_a_3_4 /= "111100110110000100010010000" OR uut_a_3_5 /= "111010111100001001010010000" OR uut_a_4_0 /= "000000000000101110100001100" OR uut_a_4_1 /= "111110001100011010101101110" OR uut_a_4_2 /= "111101000110101000011011100" OR uut_a_4_3 /= "111111111111001101100001000" OR uut_a_4_4 /= "000001111101011010110101110" OR uut_a_4_5 /= "000011001001001001001111000" OR uut_a_5_0 /= "000000000001001010100111010" OR uut_a_5_1 /= "111101000110101000011011100" OR uut_a_5_2 /= "111011010110101101100001010" OR uut_a_5_3 /= "111111111110101111000010010" OR uut_a_5_4 /= "000011001001001001001111000" OR uut_a_5_5 /= "000101000010100101110000010" THEN
              FAIL <= '1';
              FAIL_NUM <= "11000100";
              state <= "11111101";
            ELSE
              state <= "11010010";
            END IF;
            uut_rst <= '0';
          WHEN "11010010" =>
            uut_coord_shift <= "1001";
            uut_x <= "000100100011";
            uut_y <= "110111000110";
            uut_fx <= "0101011001";
            uut_fy <= "0111100010";
            uut_ft <= "0101100011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001011100110100100" OR uut_a_0_1 /= "000000011111111010000011000" OR uut_a_0_2 /= "111111010011000010100100100" OR uut_a_0_3 /= "111111111111111111001001100" OR uut_a_0_4 /= "111111111111101101010001000" OR uut_a_0_5 /= "000000000000011010011001100" OR uut_a_1_0 /= "000000000000000111111110100" OR uut_a_1_1 /= "000000000010101111011111010" OR uut_a_1_2 /= "111111111100001000101110001" OR uut_a_1_3 /= "111111111111111111111011010" OR uut_a_1_4 /= "111111111111111110011000111" OR uut_a_1_5 /= "000000000000000010010001001" OR uut_a_2_0 /= "111111111111110100110000101" OR uut_a_2_1 /= "111111111100001000101110001" OR uut_a_2_2 /= "000000000101011100011100000" OR uut_a_2_3 /= "000000000000000000000110100" OR uut_a_2_4 /= "000000000000000010010001001" OR uut_a_2_5 /= "111111111111111100110011011" OR uut_a_3_0 /= "111111111111111111001001100" OR uut_a_3_1 /= "111111111111101101010001000" OR uut_a_3_2 /= "000000000000011010011001100" OR uut_a_3_3 /= "000000000000000000000000100" OR uut_a_3_4 /= "000000000000000000001011000" OR uut_a_3_5 /= "111111111111111111110000100" OR uut_a_4_0 /= "111111111111111111111011010" OR uut_a_4_1 /= "111111111111111110011000111" OR uut_a_4_2 /= "000000000000000010010001001" OR uut_a_4_3 /= "000000000000000000000000000" OR uut_a_4_4 /= "000000000000000000000000111" OR uut_a_4_5 /= "111111111111111111111110101" OR uut_a_5_0 /= "000000000000000000000110100" OR uut_a_5_1 /= "000000000000000010010001001" OR uut_a_5_2 /= "111111111111111100110011011" OR uut_a_5_3 /= "111111111111111111111111111" OR uut_a_5_4 /= "111111111111111111111110101" OR uut_a_5_5 /= "000000000000000000000001111" THEN
              FAIL <= '1';
              FAIL_NUM <= "11000101";
              state <= "11111101";
            ELSE
              state <= "11010011";
            END IF;
            uut_rst <= '0';
          WHEN "11010011" =>
            uut_coord_shift <= "1001";
            uut_x <= "000000001100";
            uut_y <= "111000111100";
            uut_fx <= "0011111101";
            uut_fy <= "1011110011";
            uut_ft <= "0111010100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001111110000000100" OR uut_a_0_1 /= "000100000111110101000011000" OR uut_a_0_2 /= "000001001011110011010011010" OR uut_a_0_3 /= "000000000001001001111010110" OR uut_a_0_4 /= "000010011010110001000000100" OR uut_a_0_5 /= "000000101100011101110101111" OR uut_a_1_0 /= "000000000001000001111101010" OR uut_a_1_1 /= "000010001010000110010001000" OR uut_a_1_2 /= "000000100111101011010110100" OR uut_a_1_3 /= "000000000000100110101100010" OR uut_a_1_4 /= "000001010001000000101001110" OR uut_a_1_5 /= "000000010111010001100111101" OR uut_a_2_0 /= "000000000000010010111100110" OR uut_a_2_1 /= "000000100111101011010110100" OR uut_a_2_2 /= "000000001011011001100101110" OR uut_a_2_3 /= "000000000000001011000111011" OR uut_a_2_4 /= "000000010111010001100111101" OR uut_a_2_5 /= "000000000110101011111111001" OR uut_a_3_0 /= "000000000001001001111010110" OR uut_a_3_1 /= "000010011010110001000000100" OR uut_a_3_2 /= "000000101100011101110101111" OR uut_a_3_3 /= "000000000000101011010111001" OR uut_a_3_4 /= "000001011010110010011010110" OR uut_a_3_5 /= "000000011010000101011010010" OR uut_a_4_0 /= "000000000000100110101100010" OR uut_a_4_1 /= "000001010001000000101001110" OR uut_a_4_2 /= "000000010111010001100111101" OR uut_a_4_3 /= "000000000000010110101100100" OR uut_a_4_4 /= "000000101111100001011001000" OR uut_a_4_5 /= "000000001101101001110101010" OR uut_a_5_0 /= "000000000000001011000111011" OR uut_a_5_1 /= "000000010111010001100111101" OR uut_a_5_2 /= "000000000110101011111111001" OR uut_a_5_3 /= "000000000000000110100001010" OR uut_a_5_4 /= "000000001101101001110101010" OR uut_a_5_5 /= "000000000011111011000100000" THEN
              FAIL <= '1';
              FAIL_NUM <= "11000110";
              state <= "11111101";
            ELSE
              state <= "11010100";
            END IF;
            uut_rst <= '0';
          WHEN "11010100" =>
            uut_coord_shift <= "1001";
            uut_x <= "000011110110";
            uut_y <= "000011001101";
            uut_fx <= "1010110001";
            uut_fy <= "1001011101";
            uut_ft <= "1100000101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000101010101010000100" OR uut_a_0_1 /= "000000001010101010100001000" OR uut_a_0_2 /= "111001100000000101111001000" OR uut_a_0_3 /= "000000000100100110101110010" OR uut_a_0_4 /= "000000001001001101011100100" OR uut_a_0_5 /= "111010011000110011101000100" OR uut_a_1_0 /= "000000000000000010101010101" OR uut_a_1_1 /= "000000000000000101010101010" OR uut_a_1_2 /= "111111111100110000000010111" OR uut_a_1_3 /= "000000000000000010010011010" OR uut_a_1_4 /= "000000000000000100100110101" OR uut_a_1_5 /= "111111111101001100011001110" OR uut_a_2_0 /= "111111111110011000000001011" OR uut_a_2_1 /= "111111111100110000000010111" OR uut_a_2_2 /= "000001111110101110001101001" OR uut_a_2_3 /= "111111111110100110001100111" OR uut_a_2_4 /= "111111111101001100011001110" OR uut_a_2_5 /= "000001101101011100010001001" OR uut_a_3_0 /= "000000000100100110101110010" OR uut_a_3_1 /= "000000001001001101011100100" OR uut_a_3_2 /= "111010011000110011101000100" OR uut_a_3_3 /= "000000000011111110100010001" OR uut_a_3_4 /= "000000000111111101000100010" OR uut_a_3_5 /= "111011001001110010011010010" OR uut_a_4_0 /= "000000000000000010010011010" OR uut_a_4_1 /= "000000000000000100100110101" OR uut_a_4_2 /= "111111111101001100011001110" OR uut_a_4_3 /= "000000000000000001111111010" OR uut_a_4_4 /= "000000000000000011111110100" OR uut_a_4_5 /= "111111111101100100111001001" OR uut_a_5_0 /= "111111111110100110001100111" OR uut_a_5_1 /= "111111111101001100011001110" OR uut_a_5_2 /= "000001101101011100010001001" OR uut_a_5_3 /= "111111111110110010011100100" OR uut_a_5_4 /= "111111111101100100111001001" OR uut_a_5_5 /= "000001011110100001001001000" THEN
              FAIL <= '1';
              FAIL_NUM <= "11000111";
              state <= "11111101";
            ELSE
              state <= "11010101";
            END IF;
            uut_rst <= '0';
          WHEN "11010101" =>
            uut_coord_shift <= "1001";
            uut_x <= "001011011110";
            uut_y <= "001101001001";
            uut_fx <= "0011001100";
            uut_fy <= "0011100111";
            uut_ft <= "1011101011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000100110101011000" OR uut_a_0_1 /= "000001101010010110011011000" OR uut_a_0_2 /= "111111010101101100111001101" OR uut_a_0_3 /= "111111111111001111100111000" OR uut_a_0_4 /= "111101111010111011011011000" OR uut_a_0_5 /= "000000110100111011010001101" OR uut_a_1_0 /= "000000000000001101010010110" OR uut_a_1_1 /= "000000100100100011101101010" OR uut_a_1_2 /= "111111110001011101011011110" OR uut_a_1_3 /= "111111111111101111010111011" OR uut_a_1_4 /= "111111010010010000011011010" OR uut_a_1_5 /= "000000010010001100011000000" OR uut_a_2_0 /= "111111111111111010101101100" OR uut_a_2_1 /= "111111110001011101011011110" OR uut_a_2_2 /= "000000000101110010000111000" OR uut_a_2_3 /= "000000000000000110100111011" OR uut_a_2_4 /= "000000010010001100011000000" OR uut_a_2_5 /= "111111111000110000111001010" OR uut_a_3_0 /= "111111111111001111100111000" OR uut_a_3_1 /= "111101111010111011011011000" OR uut_a_3_2 /= "000000110100111011010001101" OR uut_a_3_3 /= "000000000000111100100011000" OR uut_a_3_4 /= "000010100110100000011011000" OR uut_a_3_5 /= "111110111101110001101001101" OR uut_a_4_0 /= "111111111111101111010111011" OR uut_a_4_1 /= "111111010010010000011011010" OR uut_a_4_2 /= "000000010010001100011000000" OR uut_a_4_3 /= "000000000000010100110100000" OR uut_a_4_4 /= "000000111001001111001001010" OR uut_a_4_5 /= "111111101001001111000100010" OR uut_a_5_0 /= "000000000000000110100111011" OR uut_a_5_1 /= "000000010010001100011000000" OR uut_a_5_2 /= "111111111000110000111001010" OR uut_a_5_3 /= "111111111111110111101110001" OR uut_a_5_4 /= "111111101001001111000100010" OR uut_a_5_5 /= "000000001001000011011101100" THEN
              FAIL <= '1';
              FAIL_NUM <= "11001000";
              state <= "11111101";
            ELSE
              state <= "11010110";
            END IF;
            uut_rst <= '0';
          WHEN "11010110" =>
            uut_coord_shift <= "1001";
            uut_x <= "000010011011";
            uut_y <= "001001111100";
            uut_fx <= "1110011110";
            uut_fy <= "0111110100";
            uut_ft <= "1001011100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000011001011111101000" OR uut_a_0_1 /= "000001101001001010011111000" OR uut_a_0_2 /= "110100110001011000010110011" OR uut_a_0_3 /= "000000000010111001101010000" OR uut_a_0_4 /= "000001011111101110101010000" OR uut_a_0_5 /= "110101110001110110100001000" OR uut_a_1_0 /= "000000000000001101001001010" OR uut_a_1_1 /= "000000000110110001110011010" OR uut_a_1_2 /= "111111010001101011101100011" OR uut_a_1_3 /= "000000000000001011111101110" OR uut_a_1_4 /= "000000000110001010111000011" OR uut_a_1_5 /= "111111010101110101101000111" OR uut_a_2_0 /= "111111111110100110001011000" OR uut_a_2_1 /= "111111010001101011101100011" OR uut_a_2_2 /= "000100111100100000000101101" OR uut_a_2_3 /= "111111111110101110001110110" OR uut_a_2_4 /= "111111010101110101101000111" OR uut_a_2_5 /= "000100100000000110110011010" OR uut_a_3_0 /= "000000000010111001101010000" OR uut_a_3_1 /= "000001011111101110101010000" OR uut_a_3_2 /= "110101110001110110100001000" OR uut_a_3_3 /= "000000000010101001000000000" OR uut_a_3_4 /= "000001010111001001000000000" OR uut_a_3_5 /= "110110101100100010100000000" OR uut_a_4_0 /= "000000000000001011111101110" OR uut_a_4_1 /= "000000000110001010111000011" OR uut_a_4_2 /= "111111010101110101101000111" OR uut_a_4_3 /= "000000000000001010111001001" OR uut_a_4_4 /= "000000000101100111011101001" OR uut_a_4_5 /= "111111011001100111101110010" OR uut_a_5_0 /= "111111111110101110001110110" OR uut_a_5_1 /= "111111010101110101101000111" OR uut_a_5_2 /= "000100100000000110110011010" OR uut_a_5_3 /= "111111111110110101100100010" OR uut_a_5_4 /= "111111011001100111101110010" OR uut_a_5_5 /= "000100000110010000100011100" THEN
              FAIL <= '1';
              FAIL_NUM <= "11001001";
              state <= "11111101";
            ELSE
              state <= "11010111";
            END IF;
            uut_rst <= '0';
          WHEN "11010111" =>
            uut_coord_shift <= "1001";
            uut_x <= "111010010010";
            uut_y <= "000000010111";
            uut_fx <= "1000111110";
            uut_fy <= "0011100111";
            uut_ft <= "0000111010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001110100001111000" OR uut_a_0_1 /= "110010001100011011100000000" OR uut_a_0_2 /= "000100111110101111010011011" OR uut_a_0_3 /= "000000000010100010101110101" OR uut_a_0_4 /= "101100101011000000000110100" OR uut_a_0_5 /= "000110111110001111000001101" OR uut_a_1_0 /= "111111111110010001100011011" OR uut_a_1_1 /= "001101000111100100000111100" OR uut_a_1_2 /= "111011010001001000101011010" OR uut_a_1_3 /= "111111111101100101011000000" OR uut_a_1_4 /= "010010010111011000111101110" OR uut_a_1_5 /= "111001010111111111010110001" OR uut_a_2_0 /= "000000000000100111110101111" OR uut_a_2_1 /= "111011010001001000101011010" OR uut_a_2_2 /= "000001101101010000010101101" OR uut_a_2_3 /= "000000000000110111110001111" OR uut_a_2_4 /= "111001010111111111010110001" OR uut_a_2_5 /= "000010011000111101010001101" OR uut_a_3_0 /= "000000000010100010101110101" OR uut_a_3_1 /= "101100101011000000000110100" OR uut_a_3_2 /= "000110111110001111000001101" OR uut_a_3_3 /= "000000000011100011110100100" OR uut_a_3_4 /= "100100111100001100111100010" OR uut_a_3_5 /= "001001110000101110101000101" OR uut_a_4_0 /= "111111111101100101011000000" OR uut_a_4_1 /= "010010010111011000111101110" OR uut_a_4_2 /= "111001010111111111010110001" OR uut_a_4_3 /= "111111111100100111100001100" OR uut_a_4_4 /= "011001101101100010111100111" OR uut_a_4_5 /= "110110101110011000101011111" OR uut_a_5_0 /= "000000000000110111110001111" OR uut_a_5_1 /= "111001010111111111010110001" OR uut_a_5_2 /= "000010011000111101010001101" OR uut_a_5_3 /= "000000000001001110000101110" OR uut_a_5_4 /= "110110101110011000101011111" OR uut_a_5_5 /= "000011010110001000111111000" THEN
              FAIL <= '1';
              FAIL_NUM <= "11001010";
              state <= "11111101";
            ELSE
              state <= "11011000";
            END IF;
            uut_rst <= '0';
          WHEN "11011000" =>
            uut_coord_shift <= "1001";
            uut_x <= "000000111100";
            uut_y <= "001010100011";
            uut_fx <= "0101101111";
            uut_fy <= "0100101000";
            uut_ft <= "1101000101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000100011101000000" OR uut_a_0_1 /= "111111100011111000111000110" OR uut_a_0_2 /= "000000101110110000100101010" OR uut_a_0_3 /= "000000000000101001111101111" OR uut_a_0_4 /= "111111011110111000101000001" OR uut_a_0_5 /= "000000110111000101010010110" OR uut_a_1_0 /= "111111111111111100011111000" OR uut_a_1_1 /= "000000000010110001011100111" OR uut_a_1_2 /= "111111111011011000110101010" OR uut_a_1_3 /= "111111111111111011110111000" OR uut_a_1_4 /= "000000000011010001000010100" OR uut_a_1_5 /= "111111111010100100010010100" OR uut_a_2_0 /= "000000000000000101110110000" OR uut_a_2_1 /= "111111111011011000110101010" OR uut_a_2_2 /= "000000000111101010111110000" OR uut_a_2_3 /= "000000000000000110111000101" OR uut_a_2_4 /= "111111111010100100010010100" OR uut_a_2_5 /= "000000001001000010010111100" OR uut_a_3_0 /= "000000000000101001111101111" OR uut_a_3_1 /= "111111011110111000101000001" OR uut_a_3_2 /= "000000110111000101010010110" OR uut_a_3_3 /= "000000000000110001011100000" OR uut_a_3_4 /= "111111011000111111010110110" OR uut_a_3_5 /= "000001000000111000110101010" OR uut_a_4_0 /= "111111111111111011110111000" OR uut_a_4_1 /= "000000000011010001000010100" OR uut_a_4_2 /= "111111111010100100010010100" OR uut_a_4_3 /= "111111111111111011000111111" OR uut_a_4_4 /= "000000000011110110010000000" OR uut_a_4_5 /= "111111111001100110011001001" OR uut_a_5_0 /= "000000000000000110111000101" OR uut_a_5_1 /= "111111111010100100010010100" OR uut_a_5_2 /= "000000001001000010010111100" OR uut_a_5_3 /= "000000000000001000000111000" OR uut_a_5_4 /= "111111111001100110011001001" OR uut_a_5_5 /= "000000001010101001010100101" THEN
              FAIL <= '1';
              FAIL_NUM <= "11001011";
              state <= "11111101";
            ELSE
              state <= "11011001";
            END IF;
            uut_rst <= '0';
          WHEN "11011001" =>
            uut_coord_shift <= "1001";
            uut_x <= "111110011111";
            uut_y <= "001000000100";
            uut_fx <= "1001110000";
            uut_fy <= "1001110000";
            uut_ft <= "1100010100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000110111001000" OR uut_a_0_1 /= "000000011000111110101000000" OR uut_a_0_2 /= "111111110010000111000111000" OR uut_a_0_3 /= "111111111111011111110000110" OR uut_a_0_4 /= "111110001011001000101110000" OR uut_a_0_5 /= "000001000000111110101111010" OR uut_a_1_0 /= "000000000000000011000111110" OR uut_a_1_1 /= "000000001011010100011000001" OR uut_a_1_2 /= "111111111001101101001110001" OR uut_a_1_3 /= "111111111111110001011001000" OR uut_a_1_4 /= "111111001011000010111100110" OR uut_a_1_5 /= "000000011101011100011011011" OR uut_a_2_0 /= "111111111111111110010000111" OR uut_a_2_1 /= "111111111001101101001110001" OR uut_a_2_2 /= "000000000011011111111101010" OR uut_a_2_3 /= "000000000000001000000111110" OR uut_a_2_4 /= "000000011101011100011011011" OR uut_a_2_5 /= "111111101111101000001100010" OR uut_a_3_0 /= "111111111111011111110000110" OR uut_a_3_1 /= "111110001011001000101110000" OR uut_a_3_2 /= "000001000000111110101111010" OR uut_a_3_3 /= "000000000010010110110101000" OR uut_a_3_4 /= "001000100010110000010110100" OR uut_a_3_5 /= "111011001111111111000010111" OR uut_a_4_0 /= "111111111111110001011001000" OR uut_a_4_1 /= "111111001011000010111100110" OR uut_a_4_2 /= "000000011101011100011011011" OR uut_a_4_3 /= "000000000001000100010110000" OR uut_a_4_4 /= "000011110111101111111010001" OR uut_a_4_5 /= "111101110110001111100100010" OR uut_a_5_0 /= "000000000000001000000111110" OR uut_a_5_1 /= "000000011101011100011011011" OR uut_a_5_2 /= "111111101111101000001100010" OR uut_a_5_3 /= "111111111111011001111111111" OR uut_a_5_4 /= "111101110110001111100100010" OR uut_a_5_5 /= "000001001100100110001111011" THEN
              FAIL <= '1';
              FAIL_NUM <= "11001100";
              state <= "11111101";
            ELSE
              state <= "11011010";
            END IF;
            uut_rst <= '0';
          WHEN "11011010" =>
            uut_coord_shift <= "1001";
            uut_x <= "000000110010";
            uut_y <= "001111000111";
            uut_fx <= "0011010111";
            uut_fy <= "1100111111";
            uut_ft <= "1100101010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000001001001100000" OR uut_a_0_1 /= "000001000110011111100010101" OR uut_a_0_2 /= "111111100000011010100010010" OR uut_a_0_3 /= "000000000000101100110011100" OR uut_a_0_4 /= "000101010111101111100101001" OR uut_a_0_5 /= "111101100101111110110000010" OR uut_a_1_0 /= "000000000000001000110011111" OR uut_a_1_1 /= "000001000011100110011111111" OR uut_a_1_2 /= "111111100001101101011100100" OR uut_a_1_3 /= "000000000000101010111101111" OR uut_a_1_4 /= "000101001001101001010000010" OR uut_a_1_5 /= "111101101100010011000011100" OR uut_a_2_0 /= "111111111111111100000011010" OR uut_a_2_1 /= "111111100001101101011100100" OR uut_a_2_2 /= "000000001101100100100110010" OR uut_a_2_3 /= "111111111111101100101111110" OR uut_a_2_4 /= "111101101100010011000011100" OR uut_a_2_5 /= "000001000010001011100010010" OR uut_a_3_0 /= "000000000000101100110011100" OR uut_a_3_1 /= "000101010111101111100101001" OR uut_a_3_2 /= "111101100101111110110000010" OR uut_a_3_3 /= "000000000011011010011111000" OR uut_a_3_4 /= "011010001100001100010011101" OR uut_a_3_5 /= "110100010000111101001110010" OR uut_a_4_0 /= "000000000000101010111101111" OR uut_a_4_1 /= "000101001001101001010000010" OR uut_a_4_2 /= "111101101100010011000011100" OR uut_a_4_3 /= "000000000011010001100001100" OR uut_a_4_4 /= "011001000111011100010011011" OR uut_a_4_5 /= "110100101111110000101101100" OR uut_a_5_0 /= "111111111111101100101111110" OR uut_a_5_1 /= "111101101100010011000011100" OR uut_a_5_2 /= "000001000010001011100010010" OR uut_a_5_3 /= "111111111110100010000111101" OR uut_a_5_4 /= "110100101111110000101101100" OR uut_a_5_5 /= "000101000010101101101100011" THEN
              FAIL <= '1';
              FAIL_NUM <= "11001101";
              state <= "11111101";
            ELSE
              state <= "11011011";
            END IF;
            uut_rst <= '0';
          WHEN "11011011" =>
            uut_coord_shift <= "1001";
            uut_x <= "001011001101";
            uut_y <= "001101001011";
            uut_fx <= "0010001111";
            uut_fy <= "1100000101";
            uut_ft <= "1001011011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000010111111101001100" OR uut_a_0_1 /= "110001010011101110000101011" OR uut_a_0_2 /= "111000011010111000110010111" OR uut_a_0_3 /= "111111111111001111100011000" OR uut_a_0_4 /= "000011101101101110010010000" OR uut_a_0_5 /= "000001111010101001011010000" OR uut_a_1_0 /= "111111111110001010011101110" OR uut_a_1_1 /= "001001000000101001111111001" OR uut_a_1_2 /= "000100101001100000101010110" OR uut_a_1_3 /= "000000000000011101101101110" OR uut_a_1_4 /= "111101101110001101010111011" OR uut_a_1_5 /= "111110110100110010000110110" OR uut_a_2_0 /= "111111111111000011010111000" OR uut_a_2_1 /= "000100101001100000101010110" OR uut_a_2_2 /= "000010011001011111100001111" OR uut_a_2_3 /= "000000000000001111010101001" OR uut_a_2_4 /= "111110110100110010000110110" OR uut_a_2_5 /= "111111011001001100011001100" OR uut_a_3_0 /= "111111111111001111100011000" OR uut_a_3_1 /= "000011101101101110010010000" OR uut_a_3_2 /= "000001111010101001011010000" OR uut_a_3_3 /= "000000000000001100010000000" OR uut_a_3_4 /= "111111000011111001100000000" OR uut_a_3_5 /= "111111100000111111100000000" OR uut_a_4_0 /= "000000000000011101101101110" OR uut_a_4_1 /= "111101101110001101010111011" OR uut_a_4_2 /= "111110110100110010000110110" OR uut_a_4_3 /= "111111111111111000011111001" OR uut_a_4_4 /= "000000100100110110111111001" OR uut_a_4_5 /= "000000010011000001000011101" OR uut_a_5_0 /= "000000000000001111010101001" OR uut_a_5_1 /= "111110110100110010000110110" OR uut_a_5_2 /= "111111011001001100011001100" OR uut_a_5_3 /= "111111111111111100000111111" OR uut_a_5_4 /= "000000010011000001000011101" OR uut_a_5_5 /= "000000001001110011111010001" THEN
              FAIL <= '1';
              FAIL_NUM <= "11001110";
              state <= "11111101";
            ELSE
              state <= "11011100";
            END IF;
            uut_rst <= '0';
          WHEN "11011100" =>
            uut_coord_shift <= "1010";
            uut_x <= "010101101001";
            uut_y <= "000101011011";
            uut_fx <= "0111001011";
            uut_fy <= "1000111110";
            uut_ft <= "0001010111";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000010000000000000" OR uut_a_0_1 /= "111110100111000000000000000" OR uut_a_0_2 /= "111111100101110000000000000" OR uut_a_0_3 /= "000000000000101111010000000" OR uut_a_0_4 /= "111011111001001011000000000" OR uut_a_0_5 /= "111110110010011110110000000" OR uut_a_1_0 /= "111111111111110100111000000" OR uut_a_1_1 /= "000000111101111000100000000" OR uut_a_1_2 /= "000000010010010000001000000" OR uut_a_1_3 /= "111111111111011111001001011" OR uut_a_1_4 /= "000010110110101111110110100" OR uut_a_1_5 /= "000000110101111001100111101" OR uut_a_2_0 /= "111111111111111100101110000" OR uut_a_2_1 /= "000000010010010000001000000" OR uut_a_2_2 /= "000000000101011000100010000" OR uut_a_2_3 /= "111111111111110110010011110" OR uut_a_2_4 /= "000000110101111001100111101" OR uut_a_2_5 /= "000000001111111001011100011" OR uut_a_3_0 /= "000000000000101111010000000" OR uut_a_3_1 /= "111011111001001011000000000" OR uut_a_3_2 /= "111110110010011110110000000" OR uut_a_3_3 /= "000000000010001011100010010" OR uut_a_3_4 /= "110011110111110101011111000" OR uut_a_3_5 /= "111100011011000100110011110" OR uut_a_4_0 /= "111111111111011111001001011" OR uut_a_4_1 /= "000010110110101111110110100" OR uut_a_4_2 /= "000000110101111001100111101" OR uut_a_4_3 /= "111111111110011110111110101" OR uut_a_4_4 /= "001000011011101011010011111" OR uut_a_4_5 /= "000010011111001011001010000" OR uut_a_5_0 /= "111111111111110110010011110" OR uut_a_5_1 /= "000000110101111001100111101" OR uut_a_5_2 /= "000000001111111001011100011" OR uut_a_5_3 /= "111111111111100011011000100" OR uut_a_5_4 /= "000010011111001011001010000" OR uut_a_5_5 /= "000000101110111100101000111" THEN
              FAIL <= '1';
              FAIL_NUM <= "11001111";
              state <= "11111101";
            ELSE
              state <= "11011101";
            END IF;
            uut_rst <= '0';
          WHEN "11011101" =>
            uut_coord_shift <= "1010";
            uut_x <= "110010010000";
            uut_y <= "010100111110";
            uut_fx <= "1011000100";
            uut_fy <= "1111000101";
            uut_ft <= "1110010011";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000011110101000111100" OR uut_a_0_1 /= "100110111111000100100110111" OR uut_a_0_2 /= "000111000000000110110100110" OR uut_a_0_3 /= "111111111111011011010011100" OR uut_a_0_4 /= "000011101111101010001110111" OR uut_a_0_5 /= "111110111100111010110000110" OR uut_a_1_0 /= "111111111100110111111000100" OR uut_a_1_1 /= "010100011011000000011111010" OR uut_a_1_2 /= "111010010010001010011011011" OR uut_a_1_3 /= "000000000000011101111101010" OR uut_a_1_4 /= "111100111100010101110001010" OR uut_a_1_5 /= "000000110110110001000001101" OR uut_a_2_0 /= "000000000000111000000000110" OR uut_a_2_1 /= "111010010010001010011011011" OR uut_a_2_2 /= "000001100110011001100011110" OR uut_a_2_3 /= "111111111111110111100111010" OR uut_a_2_4 /= "000000110110110001000001101" OR uut_a_2_5 /= "111111110000101010111011011" OR uut_a_3_0 /= "111111111111011011010011100" OR uut_a_3_1 /= "000011101111101010001110111" OR uut_a_3_2 /= "111110111100111010110000110" OR uut_a_3_3 /= "000000000000000101011111100" OR uut_a_3_4 /= "111111011100000111110110111" OR uut_a_3_5 /= "000000001010000010101100110" OR uut_a_4_0 /= "000000000000011101111101010" OR uut_a_4_1 /= "111100111100010101110001010" OR uut_a_4_2 /= "000000110110110001000001101" OR uut_a_4_3 /= "111111111111111011100000111" OR uut_a_4_4 /= "000000011101010010100101011" OR uut_a_4_5 /= "111111110111110011010010111" OR uut_a_5_0 /= "111111111111110111100111010" OR uut_a_5_1 /= "000000110110110001000001101" OR uut_a_5_2 /= "111111110000101010111011011" OR uut_a_5_3 /= "000000000000000001010000010" OR uut_a_5_4 /= "111111110111110011010010111" OR uut_a_5_5 /= "000000000010010010110111011" THEN
              FAIL <= '1';
              FAIL_NUM <= "11010000";
              state <= "11111101";
            ELSE
              state <= "11011110";
            END IF;
            uut_rst <= '0';
          WHEN "11011110" =>
            uut_coord_shift <= "1010";
            uut_x <= "010100111001";
            uut_y <= "001011010100";
            uut_fx <= "1011010101";
            uut_fy <= "1101000110";
            uut_ft <= "1010001001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000100111011000" OR uut_a_0_1 /= "111111101011001100010111100" OR uut_a_0_2 /= "111111111011111011000101101" OR uut_a_0_3 /= "111111111111100000110111100" OR uut_a_0_4 /= "000010000011100101001010010" OR uut_a_0_5 /= "000000011001110001111111001" OR uut_a_1_0 /= "111111111111111101011001100" OR uut_a_1_1 /= "000000001010111111100001110" OR uut_a_1_2 /= "000000000010001001110110000" OR uut_a_1_3 /= "000000000000010000011100101" OR uut_a_1_4 /= "111110111010011110111011011" OR uut_a_1_5 /= "111111110010011000010001110" OR uut_a_2_0 /= "111111111111111111011111011" OR uut_a_2_1 /= "000000000010001001110110000" OR uut_a_2_2 /= "000000000000011011000000100" OR uut_a_2_3 /= "000000000000000011001110001" OR uut_a_2_4 /= "111111110010011000010001110" OR uut_a_2_5 /= "111111111101010101001100110" OR uut_a_3_0 /= "111111111111100000110111100" OR uut_a_3_1 /= "000010000011100101001010010" OR uut_a_3_2 /= "000000011001110001111111001" OR uut_a_3_3 /= "000000000011000100111000000" OR uut_a_3_4 /= "110010111111111001000011000" OR uut_a_3_5 /= "111101011100111101100100101" OR uut_a_4_0 /= "000000000000010000011100101" OR uut_a_4_1 /= "111110111010011110111011011" OR uut_a_4_2 /= "111111110010011000010001110" OR uut_a_4_3 /= "111111111110010111111111001" OR uut_a_4_4 /= "000110110111100111101011000" OR uut_a_4_5 /= "000001010110001000101110000" OR uut_a_5_0 /= "000000000000000011001110001" OR uut_a_5_1 /= "111111110010011000010001110" OR uut_a_5_2 /= "111111111101010101001100110" OR uut_a_5_3 /= "111111111111101011100111101" OR uut_a_5_4 /= "000001010110001000101110000" OR uut_a_5_5 /= "000000010000111000001000000" THEN
              FAIL <= '1';
              FAIL_NUM <= "11010001";
              state <= "11111101";
            ELSE
              state <= "11011111";
            END IF;
            uut_rst <= '0';
          WHEN "11011111" =>
            uut_coord_shift <= "1010";
            uut_x <= "001010111110";
            uut_y <= "000100100010";
            uut_fx <= "1010101110";
            uut_fy <= "1010010111";
            uut_ft <= "1111101000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001110100001111000" OR uut_a_0_1 /= "000100001000010000001111100" OR uut_a_0_2 /= "110111111010011000111011001" OR uut_a_0_3 /= "000000000010100010011001001" OR uut_a_0_4 /= "000101110001001100000111101" OR uut_a_0_5 /= "110100101100110110000111011" OR uut_a_1_0 /= "000000000000100001000010000" OR uut_a_1_1 /= "000001001011000110000111011" OR uut_a_1_2 /= "111101101100111001111101010" OR uut_a_1_3 /= "000000000000101110001001100" OR uut_a_1_4 /= "000001101000111010101000011" OR uut_a_1_5 /= "111100110010011111101000001" OR uut_a_2_0 /= "111111111110111111010011000" OR uut_a_2_1 /= "111101101100111001111101010" OR uut_a_2_2 /= "000100100000000111111000000" OR uut_a_2_3 /= "111111111110100101100110110" OR uut_a_2_4 /= "111100110010011111101000001" OR uut_a_2_5 /= "000110010010100010011000001" OR uut_a_3_0 /= "000000000010100010011001001" OR uut_a_3_1 /= "000101110001001100000111101" OR uut_a_3_2 /= "110100101100110110000111011" OR uut_a_3_3 /= "000000000011100010111000010" OR uut_a_3_4 /= "001000000011110010111000011" OR uut_a_3_5 /= "110000001101101011100000110" OR uut_a_4_0 /= "000000000000101110001001100" OR uut_a_4_1 /= "000001101000111010101000011" OR uut_a_4_2 /= "111100110010011111101000001" OR uut_a_4_3 /= "000000000001000000011110010" OR uut_a_4_4 /= "000010010010100101000001011" OR uut_a_4_5 /= "111011100000111000110011010" OR uut_a_5_0 /= "111111111110100101100110110" OR uut_a_5_1 /= "111100110010011111101000001" OR uut_a_5_2 /= "000110010010100010011000001" OR uut_a_5_3 /= "111111111110000001101101011" OR uut_a_5_4 /= "111011100000111000110011010" OR uut_a_5_5 /= "001000110010011000101001111" THEN
              FAIL <= '1';
              FAIL_NUM <= "11010010";
              state <= "11111101";
            ELSE
              state <= "11100000";
            END IF;
            uut_rst <= '0';
          WHEN "11100000" =>
            uut_coord_shift <= "1010";
            uut_x <= "011010000111";
            uut_y <= "000011010101";
            uut_fx <= "1000100010";
            uut_fy <= "1000110111";
            uut_ft <= "0100111000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000111110100000100" OR uut_a_0_1 /= "000000000101110111000011011" OR uut_a_0_2 /= "111100100011010001000000111" OR uut_a_0_3 /= "111111111110111101100010011" OR uut_a_0_4 /= "111111111001110001001110101" OR uut_a_0_5 /= "000011101010101100011001001" OR uut_a_1_0 /= "000000000000000000101110111" OR uut_a_1_1 /= "000000000000000100011001010" OR uut_a_1_2 /= "111111111101011010011100110" OR uut_a_1_3 /= "111111111111111111001110001" OR uut_a_1_4 /= "111111111111111011010100111" OR uut_a_1_5 /= "000000000010110000000001010" OR uut_a_2_0 /= "111111111111100100011010001" OR uut_a_2_1 /= "111111111101011010011100110" OR uut_a_2_2 /= "000001100001011011101111010" OR uut_a_2_3 /= "000000000000011101010101100" OR uut_a_2_4 /= "000000000010110000000001010" OR uut_a_2_5 /= "111110011000011001111001111" OR uut_a_3_0 /= "111111111110111101100010011" OR uut_a_3_1 /= "111111111001110001001110101" OR uut_a_3_2 /= "000011101010101100011001001" OR uut_a_3_3 /= "000000000001000110101010100" OR uut_a_3_4 /= "000000000110100111111111011" OR uut_a_3_5 /= "111100000110011101101100111" OR uut_a_4_0 /= "111111111111111111001110001" OR uut_a_4_1 /= "111111111111111011010100111" OR uut_a_4_2 /= "000000000010110000000001010" OR uut_a_4_3 /= "000000000000000000110100111" OR uut_a_4_4 /= "000000000000000100111101111" OR uut_a_4_5 /= "111111111101000100110110010" OR uut_a_5_0 /= "000000000000011101010101100" OR uut_a_5_1 /= "000000000010110000000001010" OR uut_a_5_2 /= "111110011000011001111001111" OR uut_a_5_3 /= "111111111111100000110011101" OR uut_a_5_4 /= "111111111101000100110110010" OR uut_a_5_5 /= "000001101110001001011000111" THEN
              FAIL <= '1';
              FAIL_NUM <= "11010011";
              state <= "11111101";
            ELSE
              state <= "11100001";
            END IF;
            uut_rst <= '0';
          WHEN "11100001" =>
            uut_coord_shift <= "1010";
            uut_x <= "111100111001";
            uut_y <= "111000100000";
            uut_fx <= "0100101001";
            uut_fy <= "1101110101";
            uut_ft <= "0000100001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001101101100110000" OR uut_a_0_1 /= "000011010010101000001001101" OR uut_a_0_2 /= "000010101111100001011101011" OR uut_a_0_3 /= "000000000010001001000100110" OR uut_a_0_4 /= "000100000111011100001111111" OR uut_a_0_5 /= "000011011011100010001101010" OR uut_a_1_0 /= "000000000000011010010101000" OR uut_a_1_1 /= "000000110010100110011001010" OR uut_a_1_2 /= "000000101010001010101010011" OR uut_a_1_3 /= "000000000000100000111011100" OR uut_a_1_4 /= "000000111111010010011010010" OR uut_a_1_5 /= "000000110100101111010101111" OR uut_a_2_0 /= "000000000000010101111100001" OR uut_a_2_1 /= "000000101010001010101010011" OR uut_a_2_2 /= "000000100011001000111000101" OR uut_a_2_3 /= "000000000000011011011100010" OR uut_a_2_4 /= "000000110100101111010101111" OR uut_a_2_5 /= "000000101011111100110010010" OR uut_a_3_0 /= "000000000010001001000100110" OR uut_a_3_1 /= "000100000111011100001111111" OR uut_a_3_2 /= "000011011011100010001101010" OR uut_a_3_3 /= "000000000010101011011100100" OR uut_a_3_4 /= "000101001001011111111001001" OR uut_a_3_5 /= "000100010010100101001111101" OR uut_a_4_0 /= "000000000000100000111011100" OR uut_a_4_1 /= "000000111111010010011010010" OR uut_a_4_2 /= "000000110100101111010101111" OR uut_a_4_3 /= "000000000000101001001011111" OR uut_a_4_4 /= "000001001111001010000010010" OR uut_a_4_5 /= "000001000001111101101100101" OR uut_a_5_0 /= "000000000000011011011100010" OR uut_a_5_1 /= "000000110100101111010101111" OR uut_a_5_2 /= "000000101011111100110010010" OR uut_a_5_3 /= "000000000000100010010100101" OR uut_a_5_4 /= "000001000001111101101100101" OR uut_a_5_5 /= "000000110110111110000101001" THEN
              FAIL <= '1';
              FAIL_NUM <= "11010100";
              state <= "11111101";
            ELSE
              state <= "11100010";
            END IF;
            uut_rst <= '0';
          WHEN "11100010" =>
            uut_coord_shift <= "1010";
            uut_x <= "001101100010";
            uut_y <= "010111110001";
            uut_fx <= "1101010001";
            uut_fy <= "0010011010";
            uut_ft <= "0111100110";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000101000101001000" OR uut_a_0_1 /= "000011101001000011000111000" OR uut_a_0_2 /= "000100001011000001011000100" OR uut_a_0_3 /= "000000000000101110000001010" OR uut_a_0_4 /= "000100000111111001001010110" OR uut_a_0_5 /= "000100101110010111001101101" OR uut_a_1_0 /= "000000000000011101001000011" OR uut_a_1_1 /= "000010100111000011000110101" OR uut_a_1_2 /= "000010111111011001100111011" OR uut_a_1_3 /= "000000000000100000111111001" OR uut_a_1_4 /= "000010111101001010000110100" OR uut_a_1_5 /= "000011011000101110111000111" OR uut_a_2_0 /= "000000000000100001011000001" OR uut_a_2_1 /= "000010111111011001100111011" OR uut_a_2_2 /= "000011011011010011010100101" OR uut_a_2_3 /= "000000000000100101110010111" OR uut_a_2_4 /= "000011011000101110111000111" OR uut_a_2_5 /= "000011111000010100111100001" OR uut_a_3_0 /= "000000000000101110000001010" OR uut_a_3_1 /= "000100000111111001001010110" OR uut_a_3_2 /= "000100101110010111001101101" OR uut_a_3_3 /= "000000000000110100000111000" OR uut_a_3_4 /= "000100101010110100011111111" OR uut_a_3_5 /= "000101010110011000011001110" OR uut_a_4_0 /= "000000000000100000111111001" OR uut_a_4_1 /= "000010111101001010000110100" OR uut_a_4_2 /= "000011011000101110111000111" OR uut_a_4_3 /= "000000000000100101010110100" OR uut_a_4_4 /= "000011010110001100011000011" OR uut_a_4_5 /= "000011110101011010101111011" OR uut_a_5_0 /= "000000000000100101110010111" OR uut_a_5_1 /= "000011011000101110111000111" OR uut_a_5_2 /= "000011111000010100111100001" OR uut_a_5_3 /= "000000000000101010110011000" OR uut_a_5_4 /= "000011110101011010101111011" OR uut_a_5_5 /= "000100011001001100011010101" THEN
              FAIL <= '1';
              FAIL_NUM <= "11010101";
              state <= "11111101";
            ELSE
              state <= "11100011";
            END IF;
            uut_rst <= '0';
          WHEN "11100011" =>
            uut_coord_shift <= "1010";
            uut_x <= "100100111000";
            uut_y <= "000101100100";
            uut_fx <= "1110101000";
            uut_fy <= "1100111101";
            uut_ft <= "1100001110";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000001001011000010" OR uut_a_0_1 /= "000000001011010110110111011" OR uut_a_0_2 /= "000000101110100110011111100" OR uut_a_0_3 /= "111111111111010000001001100" OR uut_a_0_4 /= "111111000110000011100000010" OR uut_a_0_5 /= "111100010010001111001101000" OR uut_a_1_0 /= "000000000000000001011010110" OR uut_a_1_1 /= "000000000001101110000001100" OR uut_a_1_2 /= "000000000111000011011100111" OR uut_a_1_3 /= "111111111111111000110000011" OR uut_a_1_4 /= "111111110111001110101001111" OR uut_a_1_5 /= "111111011100000000101011010" OR uut_a_2_0 /= "000000000000000101110100110" OR uut_a_2_1 /= "000000000111000011011100111" OR uut_a_2_2 /= "000000011100111100011010000" OR uut_a_2_3 /= "111111111111100010010001111" OR uut_a_2_4 /= "111111011100000000101011010" OR uut_a_2_5 /= "111101101100010100111100010" OR uut_a_3_0 /= "111111111111010000001001100" OR uut_a_3_1 /= "111111000110000011100000010" OR uut_a_3_2 /= "111100010010001111001101000" OR uut_a_3_3 /= "000000000011110100001001000" OR uut_a_3_4 /= "000100100111101000111001100" OR uut_a_3_5 /= "010010111101000100101110000" OR uut_a_4_0 /= "111111111111111000110000011" OR uut_a_4_1 /= "111111110111001110101001111" OR uut_a_4_2 /= "111111011100000000101011010" OR uut_a_4_3 /= "000000000000100100111101000" OR uut_a_4_4 /= "000000101100110000000000001" OR uut_a_4_5 /= "000010110111100111101001101" OR uut_a_5_0 /= "111111111111100010010001111" OR uut_a_5_1 /= "111111011100000000101011010" OR uut_a_5_2 /= "111101101100010100111100010" OR uut_a_5_3 /= "000000000010010111101000100" OR uut_a_5_4 /= "000010110111100111101001101" OR uut_a_5_5 /= "001011110001011011101011100" THEN
              FAIL <= '1';
              FAIL_NUM <= "11010110";
              state <= "11111101";
            ELSE
              state <= "11100100";
            END IF;
            uut_rst <= '0';
          WHEN "11100100" =>
            uut_coord_shift <= "1010";
            uut_x <= "010000100011";
            uut_y <= "011111101100";
            uut_fx <= "1010111111";
            uut_fy <= "0100100000";
            uut_ft <= "1011001000";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000011000101110000010" OR uut_a_0_1 /= "110111001010100011000010010" OR uut_a_0_2 /= "000000100011100010001010111" OR uut_a_0_3 /= "111111111110011010011111001" OR uut_a_0_4 /= "000100100010010001000000001" OR uut_a_0_5 /= "111111101101110000100101111" OR uut_a_1_0 /= "111111111110111001010100011" OR uut_a_1_1 /= "000011001010000110101110100" OR uut_a_1_2 /= "111111110011010011001010010" OR uut_a_1_3 /= "000000000000100100010010001" OR uut_a_1_4 /= "111110011000010000001011000" OR uut_a_1_5 /= "000000000110100001010000011" OR uut_a_2_0 /= "000000000000000100011100010" OR uut_a_2_1 /= "111111110011010011001010010" OR uut_a_2_2 /= "000000000000110011000101000" OR uut_a_2_3 /= "111111111111111101101110000" OR uut_a_2_4 /= "000000000110100001010000011" OR uut_a_2_5 /= "111111111111100101110001110" OR uut_a_3_0 /= "111111111110011010011111001" OR uut_a_3_1 /= "000100100010010001000000001" OR uut_a_3_2 /= "111111101101110000100101111" OR uut_a_3_3 /= "000000000000110100000111000" OR uut_a_3_4 /= "111101101010111111110011100" OR uut_a_3_5 /= "000000001001010111010001001" OR uut_a_4_0 /= "000000000000100100010010001" OR uut_a_4_1 /= "111110011000010000001011000" OR uut_a_4_2 /= "000000000110100001010000011" OR uut_a_4_3 /= "111111111111101101010111111" OR uut_a_4_4 /= "000000110101010000011100011" OR uut_a_4_5 /= "111111111100101001110011101" OR uut_a_5_0 /= "111111111111111101101110000" OR uut_a_5_1 /= "000000000110100001010000011" OR uut_a_5_2 /= "111111111111100101110001110" OR uut_a_5_3 /= "000000000000000001001010111" OR uut_a_5_4 /= "111111111100101001110011101" OR uut_a_5_5 /= "000000000000001101011101011" THEN
              FAIL <= '1';
              FAIL_NUM <= "11010111";
              state <= "11111101";
            ELSE
              state <= "11100101";
            END IF;
            uut_rst <= '0';
          WHEN "11100101" =>
            uut_coord_shift <= "1010";
            uut_x <= "011111100000";
            uut_y <= "010011010110";
            uut_fx <= "1110110010";
            uut_fy <= "0011101010";
            uut_ft <= "1111111110";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000010000011100010000" OR uut_a_0_1 /= "000000111101101001111101111" OR uut_a_0_2 /= "001010110101101000001000000" OR uut_a_0_3 /= "000000000001101010000101100" OR uut_a_0_4 /= "000000110001101110100101000" OR uut_a_0_5 /= "001000101111011100000000010" OR uut_a_1_0 /= "000000000000000111101101001" OR uut_a_1_1 /= "000000000011100111001101011" OR uut_a_1_2 /= "000000101000101001000110011" OR uut_a_1_3 /= "000000000000000110001101110" OR uut_a_1_4 /= "000000000010111010011110101" OR uut_a_1_5 /= "000000100000110001111001000" OR uut_a_2_0 /= "000000000001010110101101000" OR uut_a_2_1 /= "000000101000101001000110011" OR uut_a_2_2 /= "000111001001001110011000110" OR uut_a_2_3 /= "000000000001000101111011100" OR uut_a_2_4 /= "000000100000110001111001000" OR uut_a_2_5 /= "000101110000110001010001011" OR uut_a_3_0 /= "000000000001101010000101100" OR uut_a_3_1 /= "000000110001101110100101000" OR uut_a_3_2 /= "001000101111011100000000010" OR uut_a_3_3 /= "000000000001010101100100000" OR uut_a_3_4 /= "000000101000000110111000000" OR uut_a_3_5 /= "000111000011001101010110000" OR uut_a_4_0 /= "000000000000000110001101110" OR uut_a_4_1 /= "000000000010111010011110101" OR uut_a_4_2 /= "000000100000110001111001000" OR uut_a_4_3 /= "000000000000000101000000110" OR uut_a_4_4 /= "000000000010010110011001110" OR uut_a_4_5 /= "000000011010011100000010000" OR uut_a_5_0 /= "000000000001000101111011100" OR uut_a_5_1 /= "000000100000110001111001000" OR uut_a_5_2 /= "000101110000110001010001011" OR uut_a_5_3 /= "000000000000111000011001101" OR uut_a_5_4 /= "000000011010011100000010000" OR uut_a_5_5 /= "000100101001011011010110111" THEN
              FAIL <= '1';
              FAIL_NUM <= "11011000";
              state <= "11111101";
            ELSE
              state <= "11100110";
            END IF;
            uut_rst <= '0';
          WHEN "11100110" =>
            uut_coord_shift <= "1010";
            uut_x <= "010011110001";
            uut_y <= "110110110101";
            uut_fx <= "1001001011";
            uut_fy <= "0001011101";
            uut_ft <= "0110100100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000010011100010000000" OR uut_a_0_1 /= "111110001001100101111000000" OR uut_a_0_2 /= "001001110101111000100000000" OR uut_a_0_3 /= "000000000010011100010000000" OR uut_a_0_4 /= "111110001001100101111000000" OR uut_a_0_5 /= "001001110101111000100000000" OR uut_a_1_0 /= "111111111111110001001100101" OR uut_a_1_1 /= "000000001011001101110110011" OR uut_a_1_2 /= "111111000100010101010101011" OR uut_a_1_3 /= "111111111111110001001100101" OR uut_a_1_4 /= "000000001011001101110110011" OR uut_a_1_5 /= "111111000100010101010101011" OR uut_a_2_0 /= "000000000001001110101111000" OR uut_a_2_1 /= "111111000100010101010101011" OR uut_a_2_2 /= "000100111101011001101110001" OR uut_a_2_3 /= "000000000001001110101111000" OR uut_a_2_4 /= "111111000100010101010101011" OR uut_a_2_5 /= "000100111101011001101110001" OR uut_a_3_0 /= "000000000010011100010000000" OR uut_a_3_1 /= "111110001001100101111000000" OR uut_a_3_2 /= "001001110101111000100000000" OR uut_a_3_3 /= "000000000010011100010000000" OR uut_a_3_4 /= "111110001001100101111000000" OR uut_a_3_5 /= "001001110101111000100000000" OR uut_a_4_0 /= "111111111111110001001100101" OR uut_a_4_1 /= "000000001011001101110110011" OR uut_a_4_2 /= "111111000100010101010101011" OR uut_a_4_3 /= "111111111111110001001100101" OR uut_a_4_4 /= "000000001011001101110110011" OR uut_a_4_5 /= "111111000100010101010101011" OR uut_a_5_0 /= "000000000001001110101111000" OR uut_a_5_1 /= "111111000100010101010101011" OR uut_a_5_2 /= "000100111101011001101110001" OR uut_a_5_3 /= "000000000001001110101111000" OR uut_a_5_4 /= "111111000100010101010101011" OR uut_a_5_5 /= "000100111101011001101110001" THEN
              FAIL <= '1';
              FAIL_NUM <= "11011001";
              state <= "11111101";
            ELSE
              state <= "11100111";
            END IF;
            uut_rst <= '0';
          WHEN "11100111" =>
            uut_coord_shift <= "1010";
            uut_x <= "101100011010";
            uut_y <= "111011101011";
            uut_fx <= "0011111111";
            uut_fy <= "1000101000";
            uut_ft <= "0111001001";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000101101001001000" OR uut_a_0_1 /= "000000010001101000100010100" OR uut_a_0_2 /= "000101010101000001111101101" OR uut_a_0_3 /= "111111111111010111011110100" OR uut_a_0_4 /= "111111110000001010111100000" OR uut_a_0_5 /= "111011001101110111011000111" OR uut_a_1_0 /= "000000000000000010001101000" OR uut_a_1_1 /= "000000000000110111000110101" OR uut_a_1_2 /= "000000010000101001101110001" OR uut_a_1_3 /= "111111111111111110000001010" OR uut_a_1_4 /= "111111111111001110100010001" OR uut_a_1_5 /= "111111110001000011010101000" OR uut_a_2_0 /= "000000000000101010101000001" OR uut_a_2_1 /= "000000010000101001101110001" OR uut_a_2_2 /= "000101000010000011000010101" OR uut_a_2_3 /= "111111111111011001101110111" OR uut_a_2_4 /= "111111110001000011010101000" OR uut_a_2_5 /= "111011011110111001111111101" OR uut_a_3_0 /= "111111111111010111011110100" OR uut_a_3_1 /= "111111110000001010111100000" OR uut_a_3_2 /= "111011001101110111011000111" OR uut_a_3_3 /= "000000000000100100011000000" OR uut_a_3_4 /= "000000001110001101011001100" OR uut_a_3_5 /= "000100010010110011110010001" OR uut_a_4_0 /= "111111111111111110000001010" OR uut_a_4_1 /= "111111111111001110100010001" OR uut_a_4_2 /= "111111110001000011010101000" OR uut_a_4_3 /= "000000000000000001110001101" OR uut_a_4_4 /= "000000000000101100011001110" OR uut_a_4_5 /= "000000001101011010110001110" OR uut_a_5_0 /= "111111111111011001101110111" OR uut_a_5_1 /= "111111110001000011010101000" OR uut_a_5_2 /= "111011011110111001111111101" OR uut_a_5_3 /= "000000000000100010010110011" OR uut_a_5_4 /= "000000001101011010110001110" OR uut_a_5_5 /= "000100000011100000110001101" THEN
              FAIL <= '1';
              FAIL_NUM <= "11011010";
              state <= "11111101";
            ELSE
              state <= "11101000";
            END IF;
            uut_rst <= '0';
          WHEN "11101000" =>
            uut_coord_shift <= "1010";
            uut_x <= "010000111000";
            uut_y <= "000011110000";
            uut_fx <= "1010111100";
            uut_fy <= "1111111110";
            uut_ft <= "0000010010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000010011111110000" OR uut_a_0_1 /= "000001101111110111001001011" OR uut_a_0_2 /= "000010000011100001001111010" OR uut_a_0_3 /= "111111111111011100111100101" OR uut_a_0_4 /= "111100111011101001111100011" OR uut_a_0_5 /= "111100011001001001101011110" OR uut_a_1_0 /= "000000000000001101111110111" OR uut_a_1_1 /= "000001001110010100110011010" OR uut_a_1_2 /= "000001011100000101101101100" OR uut_a_1_3 /= "111111111111100111011101001" OR uut_a_1_4 /= "111101110110100001010011101" OR uut_a_1_5 /= "111101011110010111000101111" OR uut_a_2_0 /= "000000000000010000011100001" OR uut_a_2_1 /= "000001011100000101101101100" OR uut_a_2_2 /= "000001101100010001011011010" OR uut_a_2_3 /= "111111111111100011001001001" OR uut_a_2_4 /= "111101011110010111000101111" OR uut_a_2_5 /= "111101000001111101001010001" OR uut_a_3_0 /= "111111111111011100111100101" OR uut_a_3_1 /= "111100111011101001111100011" OR uut_a_3_2 /= "111100011001001001101011110" OR uut_a_3_3 /= "000000000000111101100001100" OR uut_a_3_4 /= "000101011000101000100000001" OR uut_a_3_5 /= "000110010101001100100010100" OR uut_a_4_0 /= "111111111111100111011101001" OR uut_a_4_1 /= "111101110110100001010011101" OR uut_a_4_2 /= "111101011110010111000101111" OR uut_a_4_3 /= "000000000000101011000101000" OR uut_a_4_4 /= "000011110001010011110111000" OR uut_a_4_5 /= "000100011011101101110101111" OR uut_a_5_0 /= "111111111111100011001001001" OR uut_a_5_1 /= "111101011110010111000101111" OR uut_a_5_2 /= "111101000001111101001010001" OR uut_a_5_3 /= "000000000000110010101001100" OR uut_a_5_4 /= "000100011011101101110101111" OR uut_a_5_5 /= "000101001101100100110000101" THEN
              FAIL <= '1';
              FAIL_NUM <= "11011011";
              state <= "11111101";
            ELSE
              state <= "11101001";
            END IF;
            uut_rst <= '0';
          WHEN "11101001" =>
            uut_coord_shift <= "1010";
            uut_x <= "011111101000";
            uut_y <= "010110101101";
            uut_fx <= "0111011010";
            uut_fy <= "0010110111";
            uut_ft <= "1110011101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001100110110111110" OR uut_a_0_1 /= "010001011001000110100100100" OR uut_a_0_2 /= "000100010110111000001110000" OR uut_a_0_3 /= "111111111110011011001001010" OR uut_a_0_4 /= "101110111100101110010000111" OR uut_a_0_5 /= "111011101110100101101111101" OR uut_a_1_0 /= "000000000001000101100100011" OR uut_a_1_1 /= "001011110000110000011110011" OR uut_a_1_2 /= "000010111100100110001101001" OR uut_a_1_3 /= "111111111110111011110010111" OR uut_a_1_4 /= "110100011110000000001010010" OR uut_a_1_5 /= "111101000111000110011101101" OR uut_a_2_0 /= "000000000000010001011011100" OR uut_a_2_1 /= "000010111100100110001101001" OR uut_a_2_2 /= "000000101111010000000101101" OR uut_a_2_3 /= "111111111111101110111010010" OR uut_a_2_4 /= "111101000111000110011101101" OR uut_a_2_5 /= "111111010001101011001101010" OR uut_a_3_0 /= "111111111110011011001001010" OR uut_a_3_1 /= "101110111100101110010000111" OR uut_a_3_2 /= "111011101110100101101111101" OR uut_a_3_3 /= "000000000001100010111000001" OR uut_a_3_4 /= "010000101101111000010010100" OR uut_a_3_5 /= "000100001100000011001001101" OR uut_a_4_0 /= "111111111110111011110010111" OR uut_a_4_1 /= "110100011110000000001010010" OR uut_a_4_2 /= "111101000111000110011101101" OR uut_a_4_3 /= "000000000001000010110111100" OR uut_a_4_4 /= "001011010011100001101110010" OR uut_a_4_5 /= "000010110101010001100000011" OR uut_a_5_0 /= "111111111111101110111010010" OR uut_a_5_1 /= "111101000111000110011101101" OR uut_a_5_2 /= "111111010001101011001101010" OR uut_a_5_3 /= "000000000000010000110000001" OR uut_a_5_4 /= "000010110101010001100000011" OR uut_a_5_5 /= "000000101101011010101010001" THEN
              FAIL <= '1';
              FAIL_NUM <= "11011100";
              state <= "11111101";
            ELSE
              state <= "11101010";
            END IF;
            uut_rst <= '0';
          WHEN "11101010" =>
            uut_coord_shift <= "1010";
            uut_x <= "011011110101";
            uut_y <= "111110101100";
            uut_fx <= "1011101101";
            uut_fy <= "1110010110";
            uut_ft <= "0011010010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000110000110000100" OR uut_a_0_1 /= "111010110000110010100100000" OR uut_a_0_2 /= "000111111111001100011111100" OR uut_a_0_3 /= "000000000000001001000110101" OR uut_a_0_4 /= "111111000001011010011101000" OR uut_a_0_5 /= "000001011111011100011101011" OR uut_a_1_0 /= "111111111111101011000011001" OR uut_a_1_1 /= "000010010000000010010001100" OR uut_a_1_2 /= "111100100100010110001000011" OR uut_a_1_3 /= "111111111111111100000101101" OR uut_a_1_4 /= "000000011010111001001000100" OR uut_a_1_5 /= "111111010110111111010001011" OR uut_a_2_0 /= "000000000000011111111100110" OR uut_a_2_1 /= "111100100100010110001000011" OR uut_a_2_2 /= "000101001110111110001111111" OR uut_a_2_3 /= "000000000000000101111101110" OR uut_a_2_4 /= "111111010110111111010001011" OR uut_a_2_5 /= "000000111110100010101101011" OR uut_a_3_0 /= "000000000000001001000110101" OR uut_a_3_1 /= "111111000001011010011101000" OR uut_a_3_2 /= "000001011111011100011101011" OR uut_a_3_3 /= "000000000000000001101100110" OR uut_a_3_4 /= "111111110100010100001000010" OR uut_a_3_5 /= "000000010001110100100000001" OR uut_a_4_0 /= "111111111111111100000101101" OR uut_a_4_1 /= "000000011010111001001000100" OR uut_a_4_2 /= "111111010110111111010001011" OR uut_a_4_3 /= "111111111111111111010001010" OR uut_a_4_4 /= "000000000101000001010110011" OR uut_a_4_5 /= "111111111000010101111100001" OR uut_a_5_0 /= "000000000000000101111101110" OR uut_a_5_1 /= "111111010110111111010001011" OR uut_a_5_2 /= "000000111110100010101101011" OR uut_a_5_3 /= "000000000000000001000111010" OR uut_a_5_4 /= "111111111000010101111100001" OR uut_a_5_5 /= "000000001011101011010101110" THEN
              FAIL <= '1';
              FAIL_NUM <= "11011101";
              state <= "11111101";
            ELSE
              state <= "11101011";
            END IF;
            uut_rst <= '0';
          WHEN "11101011" =>
            uut_coord_shift <= "1010";
            uut_x <= "000011101111";
            uut_y <= "010000011011";
            uut_fx <= "0111111011";
            uut_fy <= "0111011010";
            uut_ft <= "0000100100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000101011101001110" OR uut_a_0_1 /= "000111000111111101111010110" OR uut_a_0_2 /= "000011110110111010010100110" OR uut_a_0_3 /= "000000000000011011001001111" OR uut_a_0_4 /= "000100011011101001010011001" OR uut_a_0_5 /= "000010011001100110001101011" OR uut_a_1_0 /= "000000000000011100011111110" OR uut_a_1_1 /= "000100101001101010111001000" OR uut_a_1_2 /= "000010100001001100010000111" OR uut_a_1_3 /= "000000000000010001101110100" OR uut_a_1_4 /= "000010111001001011000011100" OR uut_a_1_5 /= "000001100100010001011110011" OR uut_a_2_0 /= "000000000000001111011011101" OR uut_a_2_1 /= "000010100001001100010000111" OR uut_a_2_2 /= "000001010111010010010111100" OR uut_a_2_3 /= "000000000000001001100110011" OR uut_a_2_4 /= "000001100100010001011110011" OR uut_a_2_5 /= "000000110110010011001000011" OR uut_a_3_0 /= "000000000000011011001001111" OR uut_a_3_1 /= "000100011011101001010011001" OR uut_a_3_2 /= "000010011001100110001101011" OR uut_a_3_3 /= "000000000000010000111001001" OR uut_a_3_4 /= "000010110000011100101100000" OR uut_a_3_5 /= "000001011111100011000111010" OR uut_a_4_0 /= "000000000000010001101110100" OR uut_a_4_1 /= "000010111001001011000011100" OR uut_a_4_2 /= "000001100100010001011110011" OR uut_a_4_3 /= "000000000000001011000001110" OR uut_a_4_4 /= "000001110011001100001110101" OR uut_a_4_5 /= "000000111110011000001001000" OR uut_a_5_0 /= "000000000000001001100110011" OR uut_a_5_1 /= "000001100100010001011110011" OR uut_a_5_2 /= "000000110110010011001000011" OR uut_a_5_3 /= "000000000000000101111110001" OR uut_a_5_4 /= "000000111110011000001001000" OR uut_a_5_5 /= "000000100001110001110010011" THEN
              FAIL <= '1';
              FAIL_NUM <= "11011110";
              state <= "11111101";
            ELSE
              state <= "11101100";
            END IF;
            uut_rst <= '0';
          WHEN "11101100" =>
            uut_coord_shift <= "1010";
            uut_x <= "011101101100";
            uut_y <= "100111011010";
            uut_fx <= "1000110101";
            uut_fy <= "1100111000";
            uut_ft <= "0001010010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000110111110010001" OR uut_a_0_1 /= "000100110001111011111001111" OR uut_a_0_2 /= "000001111110011000100100001" OR uut_a_0_3 /= "000000000000111011100101000" OR uut_a_0_4 /= "000101000110110000010000111" OR uut_a_0_5 /= "000010000110111110111110000" OR uut_a_1_0 /= "000000000000010011000111101" OR uut_a_1_1 /= "000001101000110111011110001" OR uut_a_1_2 /= "000000101011010100100010111" OR uut_a_1_3 /= "000000000000010100011011000" OR uut_a_1_4 /= "000001110000000000001010110" OR uut_a_1_5 /= "000000101110010001001101011" OR uut_a_2_0 /= "000000000000000111111001100" OR uut_a_2_1 /= "000000101011010100100010111" OR uut_a_2_2 /= "000000010001111001010110100" OR uut_a_2_3 /= "000000000000001000011011111" OR uut_a_2_4 /= "000000101110010001001101011" OR uut_a_2_5 /= "000000010011000111010010101" OR uut_a_3_0 /= "000000000000111011100101000" OR uut_a_3_1 /= "000101000110110000010000111" OR uut_a_3_2 /= "000010000110111110111110000" OR uut_a_3_3 /= "000000000000111111101000100" OR uut_a_3_4 /= "000101011100111111010010011" OR uut_a_3_5 /= "000010010000001010110101000" OR uut_a_4_0 /= "000000000000010100011011000" OR uut_a_4_1 /= "000001110000000000001010110" OR uut_a_4_2 /= "000000101110010001001101011" OR uut_a_4_3 /= "000000000000010101110011111" OR uut_a_4_4 /= "000001110111100111111100011" OR uut_a_4_5 /= "000000110001011010101101100" OR uut_a_5_0 /= "000000000000001000011011111" OR uut_a_5_1 /= "000000101110010001001101011" OR uut_a_5_2 /= "000000010011000111010010101" OR uut_a_5_3 /= "000000000000001001000000101" OR uut_a_5_4 /= "000000110001011010101101100" OR uut_a_5_5 /= "000000010100011010100010001" THEN
              FAIL <= '1';
              FAIL_NUM <= "11011111";
              state <= "11111101";
            ELSE
              state <= "11101101";
            END IF;
            uut_rst <= '0';
          WHEN "11101101" =>
            uut_coord_shift <= "1010";
            uut_x <= "000001111110";
            uut_y <= "011001101011";
            uut_fx <= "0000101010";
            uut_fy <= "1110111010";
            uut_ft <= "0000101100";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001101111100100001" OR uut_a_0_1 /= "010110110000011100000110011" OR uut_a_0_2 /= "000010111001101001100111010" OR uut_a_0_3 /= "000000000001101010101010011" OR uut_a_0_4 /= "010101110000011101000000100" OR uut_a_0_5 /= "000010110001011111100111100" OR uut_a_1_0 /= "000000000001011011000001110" OR uut_a_1_1 /= "010010100100010101011011011" OR uut_a_1_2 /= "000010010111011110011011000" OR uut_a_1_3 /= "000000000001010111000001110" OR uut_a_1_4 /= "010001110000001000001010110" OR uut_a_1_5 /= "000010010000110100100001000" OR uut_a_2_0 /= "000000000000001011100110100" OR uut_a_2_1 /= "000010010111011110011011000" OR uut_a_2_2 /= "000000010011010011101110111" OR uut_a_2_3 /= "000000000000001011000101111" OR uut_a_2_4 /= "000010010000110100100001000" OR uut_a_2_5 /= "000000010010011101011100011" OR uut_a_3_0 /= "000000000001101010101010011" OR uut_a_3_1 /= "010101110000011101000000100" OR uut_a_3_2 /= "000010110001011111100111100" OR uut_a_3_3 /= "000000000001100101111110100" OR uut_a_3_4 /= "010100110011010001110100110" OR uut_a_3_5 /= "000010101001101100100011100" OR uut_a_4_0 /= "000000000001010111000001110" OR uut_a_4_1 /= "010001110000001000001010110" OR uut_a_4_2 /= "000010010000110100100001000" OR uut_a_4_3 /= "000000000001010011001101000" OR uut_a_4_4 /= "010000111110001101101100110" OR uut_a_4_5 /= "000010001010011101010100101" OR uut_a_5_0 /= "000000000000001011000101111" OR uut_a_5_1 /= "000010010000110100100001000" OR uut_a_5_2 /= "000000010010011101011100011" OR uut_a_5_3 /= "000000000000001010100110110" OR uut_a_5_4 /= "000010001010011101010100101" OR uut_a_5_5 /= "000000010001101001100010100" THEN
              FAIL <= '1';
              FAIL_NUM <= "11100000";
              state <= "11111101";
            ELSE
              state <= "11101110";
            END IF;
            uut_rst <= '0';
          WHEN "11101110" =>
            uut_coord_shift <= "1010";
            uut_x <= "001101100110";
            uut_y <= "100001000101";
            uut_fx <= "0100110100";
            uut_fy <= "1010010010";
            uut_ft <= "1111101010";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000101011000100100" OR uut_a_0_1 /= "111110111101000010011101001" OR uut_a_0_2 /= "111101011110011111000000100" OR uut_a_0_3 /= "111111111111101011110101111" OR uut_a_0_4 /= "000000011111010101101100010" OR uut_a_0_5 /= "000001001011100101110110100" OR uut_a_1_0 /= "111111111111111011110100001" OR uut_a_1_1 /= "000000000110100000011010101" OR uut_a_1_2 /= "000000001111101100011011001" OR uut_a_1_3 /= "000000000000000001111101010" OR uut_a_1_4 /= "111111111100111101000111000" OR uut_a_1_5 /= "111111111000101001111010100" OR uut_a_2_0 /= "111111111111110101111001111" OR uut_a_2_1 /= "000000001111101100011011001" OR uut_a_2_2 /= "000000100101110110101110111" OR uut_a_2_3 /= "000000000000000100101110010" OR uut_a_2_4 /= "111111111000101001111010100" OR uut_a_2_5 /= "111111101110010010001000001" OR uut_a_3_0 /= "111111111111101011110101111" OR uut_a_3_1 /= "000000011111010101101100010" OR uut_a_3_2 /= "000001001011100101110110100" OR uut_a_3_3 /= "000000000000001001011011110" OR uut_a_3_4 /= "111111110001010101010011110" OR uut_a_3_5 /= "111111011100100111110100100" OR uut_a_4_0 /= "000000000000000001111101010" OR uut_a_4_1 /= "111111111100111101000111000" OR uut_a_4_2 /= "111111111000101001111010100" OR uut_a_4_3 /= "111111111111111111000101010" OR uut_a_4_4 /= "000000000001011011001101011" OR uut_a_4_5 /= "000000000011011100000000010" OR uut_a_5_0 /= "000000000000000100101110010" OR uut_a_5_1 /= "111111111000101001111010100" OR uut_a_5_2 /= "111111101110010010001000001" OR uut_a_5_3 /= "111111111111111101110010011" OR uut_a_5_4 /= "000000000011011100000000010" OR uut_a_5_5 /= "000000001000010010101010101" THEN
              FAIL <= '1';
              FAIL_NUM <= "11100001";
              state <= "11111101";
            ELSE
              state <= "11101111";
            END IF;
            uut_rst <= '0';
          WHEN "11101111" =>
            uut_coord_shift <= "1010";
            uut_x <= "110000011100";
            uut_y <= "110111101000";
            uut_fx <= "0010100110";
            uut_fy <= "1010101110";
            uut_ft <= "1100011101";
            uut_valid_in <= '1';
            uut_done <= '0';
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000001110111101000" OR uut_a_0_1 /= "000001100101001010111010100" OR uut_a_0_2 /= "000010110001101100001110010" OR uut_a_0_3 /= "111111111111110010110101110" OR uut_a_0_4 /= "111110100110111110000100110" OR uut_a_0_5 /= "111101100011101000011100011" OR uut_a_1_0 /= "000000000000000110010100101" OR uut_a_1_1 /= "000000101010110001111011011" OR uut_a_1_2 /= "000001001011001000110000110" OR uut_a_1_3 /= "111111111111111010011011111" OR uut_a_1_4 /= "111111011010010110100111111" OR uut_a_1_5 /= "111110111101111000010010100" OR uut_a_2_0 /= "000000000000001011000110110" OR uut_a_2_1 /= "000001001011001000110000110" OR uut_a_2_2 /= "000010000011111101110111111" OR uut_a_2_3 /= "111111111111110110001110100" OR uut_a_2_4 /= "111110111101111000010010100" OR uut_a_2_5 /= "111110001011110111101000010" OR uut_a_3_0 /= "111111111111110010110101110" OR uut_a_3_1 /= "111110100110111110000100110" OR uut_a_3_2 /= "111101100011101000011100011" OR uut_a_3_3 /= "000000000000001011100101001" OR uut_a_3_4 /= "000001001110010110001011001" OR uut_a_3_5 /= "000010001001100110101001100" OR uut_a_4_0 /= "111111111111111010011011111" OR uut_a_4_1 /= "111111011010010110100111111" OR uut_a_4_2 /= "111110111101111000010010100" OR uut_a_4_3 /= "000000000000000100111001011" OR uut_a_4_4 /= "000000100001001000010000000" OR uut_a_4_5 /= "000000111010001011111001111" OR uut_a_5_0 /= "111111111111110110001110100" OR uut_a_5_1 /= "111110111101111000010010100" OR uut_a_5_2 /= "111110001011110111101000010" OR uut_a_5_3 /= "000000000000001000100110011" OR uut_a_5_4 /= "000000111010001011111001111" OR uut_a_5_5 /= "000001100110001100011111000" THEN
              FAIL <= '1';
              FAIL_NUM <= "11100010";
              state <= "11111101";
            ELSE
              state <= "11110000";
            END IF;
            uut_rst <= '0';
          WHEN "11110000" =>
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000011110010000" OR uut_a_0_1 /= "111111001100101101111000000" OR uut_a_0_2 /= "000000001010100001000100000" OR uut_a_0_3 /= "000000000000001000011000010" OR uut_a_0_4 /= "111110001110010111000111000" OR uut_a_0_5 /= "000000010111010011011100100" OR uut_a_1_0 /= "111111111111111100110010110" OR uut_a_1_1 /= "000000101011011110000111010" OR uut_a_1_2 /= "111111110111000101011110010" OR uut_a_1_3 /= "111111111111111000111001011" OR uut_a_1_4 /= "000001100000010100111010010" OR uut_a_1_5 /= "111111101100001111110001000" OR uut_a_2_0 /= "000000000000000000101010000" OR uut_a_2_1 /= "111111110111000101011110010" OR uut_a_2_2 /= "000000000001110100111111110" OR uut_a_2_3 /= "000000000000000001011101001" OR uut_a_2_4 /= "111111101100001111110001000" OR uut_a_2_5 /= "000000000100000011010000010" OR uut_a_3_0 /= "000000000000001000011000010" OR uut_a_3_1 /= "111110001110010111000111000" OR uut_a_3_2 /= "000000010111010011011100100" OR uut_a_3_3 /= "000000000000010010100100010" OR uut_a_3_4 /= "111100000100001011111011111" OR uut_a_3_5 /= "000000110011101000111010000" OR uut_a_4_0 /= "111111111111111000111001011" OR uut_a_4_1 /= "000001100000010100111010010" OR uut_a_4_2 /= "111111101100001111110001000" OR uut_a_4_3 /= "111111111111110000010000101" OR uut_a_4_4 /= "000011010101011100111000011" OR uut_a_4_5 /= "111111010100001110100100110" OR uut_a_5_0 /= "000000000000000001011101001" OR uut_a_5_1 /= "111111101100001111110001000" OR uut_a_5_2 /= "000000000100000011010000010" OR uut_a_5_3 /= "000000000000000011001110100" OR uut_a_5_4 /= "111111010100001110100100110" OR uut_a_5_5 /= "000000001000111110011111000" THEN
              FAIL <= '1';
              FAIL_NUM <= "11100011";
              state <= "11111101";
            ELSE
              state <= "11110001";
            END IF;
            uut_rst <= '0';
          WHEN "11110001" =>
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000110010010100000" OR uut_a_0_1 /= "000110100000010000101110100" OR uut_a_0_2 /= "001100011101001001010111101" OR uut_a_0_3 /= "111111111111010010110111000" OR uut_a_0_4 /= "111010001010100010000010100" OR uut_a_0_5 /= "110100110100110011011010000" OR uut_a_1_0 /= "000000000000011010000001000" OR uut_a_1_1 /= "000011010111001111101001100" OR uut_a_1_2 /= "000110011100001100100100000" OR uut_a_1_3 /= "111111111111101000101010001" OR uut_a_1_4 /= "111100111110111000100010011" OR uut_a_1_5 /= "111010001110001011011101001" OR uut_a_2_0 /= "000000000000110001110100100" OR uut_a_2_1 /= "000110011100001100100100000" OR uut_a_2_2 /= "001100010101010111001001110" OR uut_a_2_3 /= "111111111111010011010011001" OR uut_a_2_4 /= "111010001110001011011101001" OR uut_a_2_5 /= "110100111011110010011001110" OR uut_a_3_0 /= "111111111111010010110111000" OR uut_a_3_1 /= "111010001010100010000010100" OR uut_a_3_2 /= "110100110100110011011010000" OR uut_a_3_3 /= "000000000000101000100000000" OR uut_a_3_4 /= "000101001111000100110000000" OR uut_a_3_5 /= "001010000001101011000000000" OR uut_a_4_0 /= "111111111111101000101010001" OR uut_a_4_1 /= "111100111110111000100010011" OR uut_a_4_2 /= "111010001110001011011101001" OR uut_a_4_3 /= "000000000000010100111100010" OR uut_a_4_4 /= "000010101101010000110111001" OR uut_a_4_5 /= "000101001011110011010101000" OR uut_a_5_0 /= "111111111111010011010011001" OR uut_a_5_1 /= "111010001110001011011101001" OR uut_a_5_2 /= "110100111011110010011001110" OR uut_a_5_3 /= "000000000000101000000110101" OR uut_a_5_4 /= "000101001011110011010101000" OR uut_a_5_5 /= "001001111011011001111101001" THEN
              FAIL <= '1';
              FAIL_NUM <= "11100100";
              state <= "11111101";
            ELSE
              state <= "11110010";
            END IF;
            uut_rst <= '0';
          WHEN "11110010" =>
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000010111110001" OR uut_a_0_1 /= "000000101110110010011110000" OR uut_a_0_2 /= "000000011100101110110111011" OR uut_a_0_3 /= "111111111111110111000101101" OR uut_a_0_4 /= "111101110011101000100110000" OR uut_a_0_5 /= "111110101001110011011001111" OR uut_a_1_0 /= "000000000000000010111011001" OR uut_a_1_1 /= "000000101110000011101011100" OR uut_a_1_2 /= "000000011100010010001000100" OR uut_a_1_3 /= "111111111111110111001110100" OR uut_a_1_4 /= "111101110101110100111101011" OR uut_a_1_5 /= "111110101011001001100110011" OR uut_a_2_0 /= "000000000000000001110010111" OR uut_a_2_1 /= "000000011100010010001000100" OR uut_a_2_2 /= "000000010001010111100101000" OR uut_a_2_3 /= "111111111111111010100111001" OR uut_a_2_4 /= "111110101011001001100110011" OR uut_a_2_5 /= "111111001011111001010000101" OR uut_a_3_0 /= "111111111111110111000101101" OR uut_a_3_1 /= "111101110011101000100110000" OR uut_a_3_2 /= "111110101001110011011001111" OR uut_a_3_3 /= "000000000000011010101111001" OR uut_a_3_4 /= "000110100101000110001110000" OR uut_a_3_5 /= "000100000010100101110010011" OR uut_a_4_0 /= "111111111111110111001110100" OR uut_a_4_1 /= "111101110101110100111101011" OR uut_a_4_2 /= "111110101011001001100110011" OR uut_a_4_3 /= "000000000000011010010100011" OR uut_a_4_4 /= "000110011110100001000111110" OR uut_a_4_5 /= "000011111110100011001100100" OR uut_a_5_0 /= "111111111111111010100111001" OR uut_a_5_1 /= "111110101011001001100110011" OR uut_a_5_2 /= "111111001011111001010000101" OR uut_a_5_3 /= "000000000000010000001010010" OR uut_a_5_4 /= "000011111110100011001100100" OR uut_a_5_5 /= "000010011100010100001101111" THEN
              FAIL <= '1';
              FAIL_NUM <= "11100101";
              state <= "11111101";
            ELSE
              state <= "11110011";
            END IF;
            uut_rst <= '0';
          WHEN "11110011" =>
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001011101001111110" OR uut_a_0_1 /= "001110011001100010011101101" OR uut_a_0_2 /= "111001010100011000001000001" OR uut_a_0_3 /= "111111111111101100001001111" OR uut_a_0_4 /= "111100111011111000100001001" OR uut_a_0_5 /= "000001011011000000010010001" OR uut_a_1_0 /= "000000000000111001100110001" OR uut_a_1_1 /= "001000111001001101100100010" OR uut_a_1_2 /= "111011110111110111100001110" OR uut_a_1_3 /= "111111111111110011101111100" OR uut_a_1_4 /= "111110000110110111010000010" OR uut_a_1_5 /= "000000111000001101100001001" OR uut_a_2_0 /= "111111111111100101010001100" OR uut_a_2_1 /= "111011110111110111100001110" OR uut_a_2_2 /= "000001111010100100001101011" OR uut_a_2_3 /= "000000000000000101101100000" OR uut_a_2_4 /= "000000111000001101100001001" OR uut_a_2_5 /= "111111100101111010101000110" OR uut_a_3_0 /= "111111111111101100001001111" OR uut_a_3_1 /= "111100111011111000100001001" OR uut_a_3_2 /= "000001011011000000010010001" OR uut_a_3_3 /= "000000000000000100001110010" OR uut_a_3_4 /= "000000101001101111001000111" OR uut_a_3_5 /= "111111101100101000100000011" OR uut_a_4_0 /= "111111111111110011101111100" OR uut_a_4_1 /= "111110000110110111010000010" OR uut_a_4_2 /= "000000111000001101100001001" OR uut_a_4_3 /= "000000000000000010100110111" OR uut_a_4_4 /= "000000011001110001111001011" OR uut_a_4_5 /= "111111110100000010011001010" OR uut_a_5_0 /= "000000000000000101101100000" OR uut_a_5_1 /= "000000111000001101100001001" OR uut_a_5_2 /= "111111100101111010101000110" OR uut_a_5_3 /= "111111111111111110110010100" OR uut_a_5_4 /= "111111110100000010011001010" OR uut_a_5_5 /= "000000000101100011010000111" THEN
              FAIL <= '1';
              FAIL_NUM <= "11100110";
              state <= "11111101";
            ELSE
              state <= "11110100";
            END IF;
            uut_rst <= '0';
          WHEN "11110100" =>
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000011111110000000" OR uut_a_0_1 /= "111011001000111100011100011" OR uut_a_0_2 /= "111110111011010010100011101" OR uut_a_0_3 /= "111111111111000101001110110" OR uut_a_0_4 /= "001000111111110000011111110" OR uut_a_0_5 /= "000001111111001011100101001" OR uut_a_1_0 /= "111111111111101100100011110" OR uut_a_1_1 /= "000010111110011101011111010" OR uut_a_1_2 /= "000000101010000100100100110" OR uut_a_1_3 /= "000000000000100011111111000" OR uut_a_1_4 /= "111010011111011101011111100" OR uut_a_1_5 /= "111110110010001000000110001" OR uut_a_2_0 /= "111111111111111011101101001" OR uut_a_2_1 /= "000000101010000100100100110" OR uut_a_2_2 /= "000000001001010010110001010" OR uut_a_2_3 /= "000000000000000111111100101" OR uut_a_2_4 /= "111110110010001000000110001" OR uut_a_2_5 /= "111111101110110011000101110" OR uut_a_3_0 /= "111111111111000101001110110" OR uut_a_3_1 /= "001000111111110000011111110" OR uut_a_3_2 /= "000001111111001011100101001" OR uut_a_3_3 /= "000000000001101100110010000" OR uut_a_3_4 /= "101111010110010010001010000" OR uut_a_3_5 /= "111100010100100101110011000" OR uut_a_4_0 /= "000000000000100011111111000" OR uut_a_4_1 /= "111010011111011101011111100" OR uut_a_4_2 /= "111110110010001000000110001" OR uut_a_4_3 /= "111111111110111101011001001" OR uut_a_4_4 /= "001010001100100010110000100" OR uut_a_4_5 /= "000010010000001001000110110" OR uut_a_5_0 /= "000000000000000111111100101" OR uut_a_5_1 /= "111110110010001000000110001" OR uut_a_5_2 /= "111111101110110011000101110" OR uut_a_5_3 /= "111111111111110001010010010" OR uut_a_5_4 /= "000010010000001001000110110" OR uut_a_5_5 /= "000000011111110101110000110" THEN
              FAIL <= '1';
              FAIL_NUM <= "11100111";
              state <= "11111101";
            ELSE
              state <= "11110101";
            END IF;
            uut_rst <= '0';
          WHEN "11110101" =>
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000110011010000100" OR uut_a_0_1 /= "000110110000011111001110000" OR uut_a_0_2 /= "000001100000000110111100000" OR uut_a_0_3 /= "000000000000000000010100010" OR uut_a_0_4 /= "000000000010101010110111000" OR uut_a_0_5 /= "000000000000100101111110000" OR uut_a_1_0 /= "000000000000011011000001111" OR uut_a_1_1 /= "000011100100000100011101101" OR uut_a_1_2 /= "000000110010101011101010001" OR uut_a_1_3 /= "000000000000000000001010101" OR uut_a_1_4 /= "000000000001011010000110100" OR uut_a_1_5 /= "000000000000010100000001011" OR uut_a_2_0 /= "000000000000000110000000011" OR uut_a_2_1 /= "000000110010101011101010001" OR uut_a_2_2 /= "000000001011010000110100000" OR uut_a_2_3 /= "000000000000000000000010010" OR uut_a_2_4 /= "000000000000010100000001011" OR uut_a_2_5 /= "000000000000000100011100110" OR uut_a_3_0 /= "000000000000000000010100010" OR uut_a_3_1 /= "000000000010101010110111000" OR uut_a_3_2 /= "000000000000100101111110000" OR uut_a_3_3 /= "000000000000000000000000001" OR uut_a_3_4 /= "000000000000000001000011100" OR uut_a_3_5 /= "000000000000000000001111000" OR uut_a_4_0 /= "000000000000000000001010101" OR uut_a_4_1 /= "000000000001011010000110100" OR uut_a_4_2 /= "000000000000010100000001011" OR uut_a_4_3 /= "000000000000000000000000000" OR uut_a_4_4 /= "000000000000000000100011100" OR uut_a_4_5 /= "000000000000000000000111111" OR uut_a_5_0 /= "000000000000000000000010010" OR uut_a_5_1 /= "000000000000010100000001011" OR uut_a_5_2 /= "000000000000000100011100110" OR uut_a_5_3 /= "000000000000000000000000000" OR uut_a_5_4 /= "000000000000000000000111111" OR uut_a_5_5 /= "000000000000000000000001110" THEN
              FAIL <= '1';
              FAIL_NUM <= "11101000";
              state <= "11111101";
            ELSE
              state <= "11110110";
            END IF;
            uut_rst <= '0';
          WHEN "11110110" =>
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001101101101101001" OR uut_a_0_1 /= "011011000110101101100010100" OR uut_a_0_2 /= "010011011101010100101111010" OR uut_a_0_3 /= "000000000000101010010110101" OR uut_a_0_4 /= "001010011101101110101111110" OR uut_a_0_5 /= "000111100000110010100010011" OR uut_a_1_0 /= "000000000001101100011010110" OR uut_a_1_1 /= "011010110010011000100000010" OR uut_a_1_2 /= "010011001110101110101111110" OR uut_a_1_3 /= "000000000000101001110110111" OR uut_a_1_4 /= "001010010101111000011100101" OR uut_a_1_5 /= "000111011011001001111100100" OR uut_a_2_0 /= "000000000001001101110101010" OR uut_a_2_1 /= "010011001110101110101111110" OR uut_a_2_2 /= "001101110011100001011111101" OR uut_a_2_3 /= "000000000000011110000011001" OR uut_a_2_4 /= "000111011011001001111100100" OR uut_a_2_5 /= "000101010101000110110110110" OR uut_a_3_0 /= "000000000000101010010110101" OR uut_a_3_1 /= "001010011101101110101111110" OR uut_a_3_2 /= "000111100000110010100010011" OR uut_a_3_3 /= "000000000000010000010110100" OR uut_a_3_4 /= "000100000010100100010001101" OR uut_a_3_5 /= "000010111001100111110000111" OR uut_a_4_0 /= "000000000000101001110110111" OR uut_a_4_1 /= "001010010101111000011100101" OR uut_a_4_2 /= "000111011011001001111100100" OR uut_a_4_3 /= "000000000000010000001010010" OR uut_a_4_4 /= "000011111111100010010110011" OR uut_a_4_5 /= "000010110111011100100011001" OR uut_a_5_0 /= "000000000000011110000011001" OR uut_a_5_1 /= "000111011011001001111100100" OR uut_a_5_2 /= "000101010101000110110110110" OR uut_a_5_3 /= "000000000000001011100110011" OR uut_a_5_4 /= "000010110111011100100011001" OR uut_a_5_5 /= "000010000011101100010111100" THEN
              FAIL <= '1';
              FAIL_NUM <= "11101001";
              state <= "11111101";
            ELSE
              state <= "11110111";
            END IF;
            uut_rst <= '0';
          WHEN "11110111" =>
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000100100111011010" OR uut_a_0_1 /= "001000000001110010110101111" OR uut_a_0_2 /= "111111100111110001000110001" OR uut_a_0_3 /= "000000000000001110001110111" OR uut_a_0_4 /= "000011000110000010110101110" OR uut_a_0_5 /= "111111110110101010001100101" OR uut_a_1_0 /= "000000000000100000000111001" OR uut_a_1_1 /= "000110111110110011110111101" OR uut_a_1_2 /= "111111101010111011010010100" OR uut_a_1_3 /= "000000000000001100011000001" OR uut_a_1_4 /= "000010101100001110011010001" OR uut_a_1_5 /= "111111110111111000001000100" OR uut_a_2_0 /= "111111111111111110011111000" OR uut_a_2_1 /= "111111101010111011010010100" OR uut_a_2_2 /= "000000000000111111100111000" OR uut_a_2_3 /= "111111111111111111011010101" OR uut_a_2_4 /= "111111110111111000001000100" OR uut_a_2_5 /= "000000000000011000100001001" OR uut_a_3_0 /= "000000000000001110001110111" OR uut_a_3_1 /= "000011000110000010110101110" OR uut_a_3_2 /= "111111110110101010001100101" OR uut_a_3_3 /= "000000000000000101011111001" OR uut_a_3_4 /= "000001001100010101100100110" OR uut_a_3_5 /= "111111111100011001100100110" OR uut_a_4_0 /= "000000000000001100011000001" OR uut_a_4_1 /= "000010101100001110011010001" OR uut_a_4_2 /= "111111110111111000001000100" OR uut_a_4_3 /= "000000000000000100110001010" OR uut_a_4_4 /= "000001000010011000101000110" OR uut_a_4_5 /= "111111111100110111100111010" OR uut_a_5_0 /= "111111111111111111011010101" OR uut_a_5_1 /= "111111110111111000001000100" OR uut_a_5_2 /= "000000000000011000100001001" OR uut_a_5_3 /= "111111111111111111110001100" OR uut_a_5_4 /= "111111111100110111100111010" OR uut_a_5_5 /= "000000000000001001011100110" THEN
              FAIL <= '1';
              FAIL_NUM <= "11101010";
              state <= "11111101";
            ELSE
              state <= "11111000";
            END IF;
            uut_rst <= '0';
          WHEN "11111000" =>
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001111101100000110" OR uut_a_0_1 /= "000011101010010110101101010" OR uut_a_0_2 /= "010000000110100100101010100" OR uut_a_0_3 /= "000000000001110101010101111" OR uut_a_0_4 /= "000011011011000110011101100" OR uut_a_0_5 /= "001111000011011111101000001" OR uut_a_1_0 /= "000000000000001110101001011" OR uut_a_1_1 /= "000000011011010110010101100" OR uut_a_1_2 /= "000001111000010001000101110" OR uut_a_1_3 /= "000000000000001101101100011" OR uut_a_1_4 /= "000000011001100100011010010" OR uut_a_1_5 /= "000001110000011100000110001" OR uut_a_2_0 /= "000000000001000000011010010" OR uut_a_2_1 /= "000001111000010001000101110" OR uut_a_2_2 /= "001000010000110111111000001" OR uut_a_2_3 /= "000000000000111100001101111" OR uut_a_2_4 /= "000001110000011100000110001" OR uut_a_2_5 /= "000111101110011100110000110" OR uut_a_3_0 /= "000000000001110101010101111" OR uut_a_3_1 /= "000011011011000110011101100" OR uut_a_3_2 /= "001111000011011111101000001" OR uut_a_3_3 /= "000000000001101101101101001" OR uut_a_3_4 /= "000011001100110101110000011" OR uut_a_3_5 /= "001110000100110010000001001" OR uut_a_4_0 /= "000000000000001101101100011" OR uut_a_4_1 /= "000000011001100100011010010" OR uut_a_4_2 /= "000001110000011100000110001" OR uut_a_4_3 /= "000000000000001100110011010" OR uut_a_4_4 /= "000000010111111001111001011" OR uut_a_4_5 /= "000001101001000111101101100" OR uut_a_5_0 /= "000000000000111100001101111" OR uut_a_5_1 /= "000001110000011100000110001" OR uut_a_5_2 /= "000111101110011100110000110" OR uut_a_5_3 /= "000000000000111000010011001" OR uut_a_5_4 /= "000001101001000111101101100" OR uut_a_5_5 /= "000111001110010001000010110" THEN
              FAIL <= '1';
              FAIL_NUM <= "11101011";
              state <= "11111101";
            ELSE
              state <= "11111001";
            END IF;
            uut_rst <= '0';
          WHEN "11111001" =>
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000001100110110111110" OR uut_a_0_1 /= "010111110111000000000000001" OR uut_a_0_2 /= "101100001111000000000100001" OR uut_a_0_3 /= "000000000000101100110100110" OR uut_a_0_4 /= "001010011001010111000000100" OR uut_a_0_5 /= "110111011000110011010101110" OR uut_a_1_0 /= "000000000001011111011100000" OR uut_a_1_1 /= "010110001000101001101000001" OR uut_a_1_2 /= "101101101010011010101011110" OR uut_a_1_3 /= "000000000000101001100101011" OR uut_a_1_4 /= "001001101001010001101110000" OR uut_a_1_5 /= "111000000000101000101000010" OR uut_a_2_0 /= "111111111110110000111100000" OR uut_a_2_1 /= "101101101010011010101011110" OR uut_a_2_2 /= "001111001100001110001000110" OR uut_a_2_3 /= "111111111111011101100011001" OR uut_a_2_4 /= "111000000000101000101000010" OR uut_a_2_5 /= "000110100111101000000010101" OR uut_a_3_0 /= "000000000000101100110100110" OR uut_a_3_1 /= "001010011001010111000000100" OR uut_a_3_2 /= "110111011000110011010101110" OR uut_a_3_3 /= "000000000000010011100010000" OR uut_a_3_4 /= "000100100001111010101100000" OR uut_a_3_5 /= "111100001111110100111010000" OR uut_a_4_0 /= "000000000000101001100101011" OR uut_a_4_1 /= "001001101001010001101110000" OR uut_a_4_2 /= "111000000000101000101000010" OR uut_a_4_3 /= "000000000000010010000111101" OR uut_a_4_4 /= "000100001100111101110100100" OR uut_a_4_5 /= "111100100001001011101101010" OR uut_a_5_0 /= "111111111111011101100011001" OR uut_a_5_1 /= "111000000000101000101000010" OR uut_a_5_2 /= "000110100111101000000010101" OR uut_a_5_3 /= "111111111111110000111111010" OR uut_a_5_4 /= "111100100001001011101101010" OR uut_a_5_5 /= "000010111000100101100001101" THEN
              FAIL <= '1';
              FAIL_NUM <= "11101100";
              state <= "11111101";
            ELSE
              state <= "11111010";
            END IF;
            uut_rst <= '0';
          WHEN "11111010" =>
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000000000110111001" OR uut_a_0_1 /= "000000000000110110010000111" OR uut_a_0_2 /= "000000001011000011100101001" OR uut_a_0_3 /= "111111111111111110100100001" OR uut_a_0_4 /= "111111111110100101100011111" OR uut_a_0_5 /= "111111101101100100101100101" OR uut_a_1_0 /= "000000000000000000000011011" OR uut_a_1_1 /= "000000000000000011010101101" OR uut_a_1_2 /= "000000000000101011100010000" OR uut_a_1_3 /= "111111111111111111111010010" OR uut_a_1_4 /= "111111111111111010011011111" OR uut_a_1_5 /= "111111111110110111011100011" OR uut_a_2_0 /= "000000000000000000101100001" OR uut_a_2_1 /= "000000000000101011100010000" OR uut_a_2_2 /= "000000001000110111101001110" OR uut_a_2_3 /= "111111111111111110110110010" OR uut_a_2_4 /= "111111111110110111011100011" OR uut_a_2_5 /= "111111110001001101111010001" OR uut_a_3_0 /= "111111111111111110100100001" OR uut_a_3_1 /= "111111111110100101100011111" OR uut_a_3_2 /= "111111101101100100101100101" OR uut_a_3_3 /= "000000000000000010011001001" OR uut_a_3_4 /= "000000000010010110101110111" OR uut_a_3_5 /= "000000011110101101100000001" OR uut_a_4_0 /= "111111111111111111111010010" OR uut_a_4_1 /= "111111111111111010011011111" OR uut_a_4_2 /= "111111111110110111011100011" OR uut_a_4_3 /= "000000000000000000001001011" OR uut_a_4_4 /= "000000000000001001010001100" OR uut_a_4_5 /= "000000000001111000111011001" OR uut_a_5_0 /= "111111111111111110110110010" OR uut_a_5_1 /= "111111111110110111011100011" OR uut_a_5_2 /= "111111110001001101111010001" OR uut_a_5_3 /= "000000000000000001111010110" OR uut_a_5_4 /= "000000000001111000111011001" OR uut_a_5_5 /= "000000011000101000110100010" THEN
              FAIL <= '1';
              FAIL_NUM <= "11101101";
              state <= "11111101";
            ELSE
              state <= "11111011";
            END IF;
            uut_rst <= '0';
          WHEN "11111011" =>
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000101110010100100" OR uut_a_0_1 /= "000100111010110101010101100" OR uut_a_0_2 /= "110100110011110110000011010" OR uut_a_0_3 /= "111111111111001000111101010" OR uut_a_0_4 /= "111010001001111000010011110" OR uut_a_0_5 /= "001101010011000001000001001" OR uut_a_1_0 /= "000000000000010011101011010" OR uut_a_1_1 /= "000010000101101111100010000" OR uut_a_1_2 /= "111011001111110001100001100" OR uut_a_1_3 /= "111111111111101000100111100" OR uut_a_1_4 /= "111101100001000100100110111" OR uut_a_1_5 /= "000101101001100000111111101" OR uut_a_2_0 /= "111111111111010011001111011" OR uut_a_2_1 /= "111011001111110001100001100" OR uut_a_2_2 /= "001010110100000001101111010" OR uut_a_2_3 /= "000000000000110101001100000" OR uut_a_2_4 /= "000101101001100000111111101" OR uut_a_2_5 /= "110011001001101001111111000" OR uut_a_3_0 /= "111111111111001000111101010" OR uut_a_3_1 /= "111010001001111000010011110" OR uut_a_3_2 /= "001101010011000001000001001" OR uut_a_3_3 /= "000000000001000001011010001" OR uut_a_3_4 /= "000110111100100100100100011" OR uut_a_3_5 /= "110000001100101110100101010" OR uut_a_4_0 /= "111111111111101000100111100" OR uut_a_4_1 /= "111101100001000100100110111" OR uut_a_4_2 /= "000101101001100000111111101" OR uut_a_4_3 /= "000000000000011011110010010" OR uut_a_4_4 /= "000010111100110110110010001" OR uut_a_4_5 /= "111001010010011010000010011" OR uut_a_5_0 /= "000000000000110101001100000" OR uut_a_5_1 /= "000101101001100000111111101" OR uut_a_5_2 /= "110011001001101001111111000" OR uut_a_5_3 /= "111111111111000000110010111" OR uut_a_5_4 /= "111001010010011010000010011" OR uut_a_5_5 /= "001111010001001100110111001" THEN
              FAIL <= '1';
              FAIL_NUM <= "11101110";
              state <= "11111101";
            ELSE
              state <= "11111100";
            END IF;
            uut_rst <= '0';
          WHEN "11111100" =>
            IF uut_valid_out /= '1' OR uut_done_buf /= '0' OR uut_a_0_0 /= "000000000000001101011101001" OR uut_a_0_1 /= "111110010111010011010111110" OR uut_a_0_2 /= "111111000111101010000010100" OR uut_a_0_3 /= "111111111111100100100110101" OR uut_a_0_4 /= "000011010101001011011100110" OR uut_a_0_5 /= "000001110010101110010000100" OR uut_a_1_0 /= "111111111111111001011101001" OR uut_a_1_1 /= "000000110010111010101101000" OR uut_a_1_2 /= "000000011011011001101011100" OR uut_a_1_3 /= "000000000000001101010100101" OR uut_a_1_4 /= "111110011000010100110011101" OR uut_a_1_5 /= "111111001000001101010000001" OR uut_a_2_0 /= "111111111111111100011110101" OR uut_a_2_1 /= "000000011011011001101011100" OR uut_a_2_2 /= "000000001110101111101111110" OR uut_a_2_3 /= "000000000000000111001010111" OR uut_a_2_4 /= "111111001000001101010000001" OR uut_a_2_5 /= "111111100001111110011001001" OR uut_a_3_0 /= "111111111111100100100110101" OR uut_a_3_1 /= "000011010101001011011100110" OR uut_a_3_2 /= "000001110010101110010000100" OR uut_a_3_3 /= "000000000000110111110010001" OR uut_a_3_4 /= "111001001101111011111101110" OR uut_a_3_5 /= "111100010110011010000110100" OR uut_a_4_0 /= "000000000000001101010100101" OR uut_a_4_1 /= "111110011000010100110011101" OR uut_a_4_2 /= "111111001000001101010000001" OR uut_a_4_3 /= "111111111111100100110111101" OR uut_a_4_4 /= "000011010011000110001101100" OR uut_a_4_5 /= "000001110001100110100011100" OR uut_a_5_0 /= "000000000000000111001010111" OR uut_a_5_1 /= "111111001000001101010000001" OR uut_a_5_2 /= "111111100001111110011001001" OR uut_a_5_3 /= "111111111111110001011001101" OR uut_a_5_4 /= "000001110001100110100011100" OR uut_a_5_5 /= "000000111101001000101010110" THEN
              FAIL <= '1';
              FAIL_NUM <= "11101111";
              state <= "11111101";
            ELSE
              state <= "11111101";
            END IF;
            uut_rst <= '0';
          WHEN OTHERS =>
            DONE <= '1';
            uut_rst <= '1';
        END CASE;
      END IF;
    END IF;
  END PROCESS;
END;
