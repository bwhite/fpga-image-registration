LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
ENTITY unscale_h_matrixT0_tb IS
PORT(
  CLK : IN STD_LOGIC;
  RST : IN STD_LOGIC;
  DONE : OUT STD_LOGIC;
  FAIL : OUT STD_LOGIC;
  FAIL_NUM : OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END unscale_h_matrixT0_tb;
ARCHITECTURE behavior OF unscale_h_matrixT0_tb IS
  COMPONENT unscale_h_matrix
  PORT(
    CLK : IN STD_LOGIC;
    RST : IN STD_LOGIC;
    H_0_0_I : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    H_0_1_I : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    H_0_2_I : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    H_1_0_I : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    H_1_1_I : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    H_1_2_I : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    XB : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    YB : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    INPUT_VALID : IN STD_LOGIC;
    H_0_0 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    H_0_1 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    H_0_2 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    H_1_0 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    H_1_1 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    H_1_2 : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    OUTPUT_VALID : OUT STD_LOGIC);
  END COMPONENT;
  SIGNAL uut_rst_wire, uut_rst : STD_LOGIC;
  SIGNAL state : STD_LOGIC_VECTOR(6 DOWNTO 0);
  -- UUT Input
  SIGNAL uut_input_valid : STD_LOGIC;
  SIGNAL uut_h_0_0_i, uut_h_0_1_i, uut_h_0_2_i, uut_h_1_0_i, uut_h_1_1_i, uut_h_1_2_i, uut_xb, uut_yb : STD_LOGIC_VECTOR(26 DOWNTO 0);
  -- UUT Output
  SIGNAL uut_output_valid : STD_LOGIC;
  SIGNAL uut_h_0_0, uut_h_0_1, uut_h_0_2, uut_h_1_0, uut_h_1_1, uut_h_1_2 : STD_LOGIC_VECTOR(26 DOWNTO 0);
BEGIN
  uut_rst_wire <= RST OR uut_rst;
  uut :  unscale_h_matrix PORT MAP (
    CLK => CLK,
    RST => uut_rst_wire,
    H_0_0_I => uut_h_0_0_i,
    H_0_1_I => uut_h_0_1_i,
    H_0_2_I => uut_h_0_2_i,
    H_1_0_I => uut_h_1_0_i,
    H_1_1_I => uut_h_1_1_i,
    H_1_2_I => uut_h_1_2_i,
    XB => uut_xb,
    YB => uut_yb,
    INPUT_VALID => uut_input_valid,
    H_0_0 => uut_h_0_0,
    H_0_1 => uut_h_0_1,
    H_0_2 => uut_h_0_2,
    H_1_0 => uut_h_1_0,
    H_1_1 => uut_h_1_1,
    H_1_2 => uut_h_1_2,
    OUTPUT_VALID => uut_output_valid
  );
  PROCESS (CLK) IS
  BEGIN
    IF CLK'event AND CLK='1' THEN
      IF RST='1' THEN
        DONE <= '0';
        FAIL <= '0';
        uut_rst <= '1';
        FAIL_NUM <= (OTHERS => '0');
        state <= (OTHERS => '0');
      ELSE
        CASE state IS
          WHEN "0000000" =>
            uut_h_0_0_i <= "111111111000010010011001010";
            uut_h_0_1_i <= "000000000101001001001011011";
            uut_h_0_2_i <= "111111110000011010101000011";
            uut_h_1_0_i <= "111111110001011101111110001";
            uut_h_1_1_i <= "111111111010100010101000011";
            uut_h_1_2_i <= "000000000110111110100110100";
            uut_xb <= "111111110001000100100111100";
            uut_yb <= "111111111100111111100001010";
            uut_input_valid <= '1';
            state <= "0000001";
            uut_rst <= '0';
          WHEN "0000001" =>
            uut_h_0_0_i <= "000000000110111010111111110";
            uut_h_0_1_i <= "000000001111011110000010111";
            uut_h_0_2_i <= "000000001001101000010111100";
            uut_h_1_0_i <= "000000001101011110111001011";
            uut_h_1_1_i <= "000000001100101011101000101";
            uut_h_1_2_i <= "000000000001110000100110001";
            uut_xb <= "111111110100000100010110001";
            uut_yb <= "000000000100111100101010011";
            uut_input_valid <= '1';
            state <= "0000010";
            uut_rst <= '0';
          WHEN "0000010" =>
            uut_h_0_0_i <= "000000001011101001011001100";
            uut_h_0_1_i <= "111111110010010000111010000";
            uut_h_0_2_i <= "111111110100111001001011101";
            uut_h_1_0_i <= "111111111000110010011000001";
            uut_h_1_1_i <= "111111111100000111110001000";
            uut_h_1_2_i <= "000000000100001100010010011";
            uut_xb <= "000000001110101100010000101";
            uut_yb <= "111111111111111101010010001";
            uut_input_valid <= '1';
            state <= "0000011";
            uut_rst <= '0';
          WHEN "0000011" =>
            uut_h_0_0_i <= "000000000111101000101010111";
            uut_h_0_1_i <= "000000000010011100100100101";
            uut_h_0_2_i <= "000000001100000110100111001";
            uut_h_1_0_i <= "111111110000011010000111111";
            uut_h_1_1_i <= "000000001001110101100000110";
            uut_h_1_2_i <= "000000001100111000000011110";
            uut_xb <= "111111110110001010011001110";
            uut_yb <= "000000001001010011111010110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111000010010011001010" OR uut_h_0_1 /= "000000000101001001001011011" OR uut_h_0_2 /= "111111011011010000100110001" OR uut_h_1_0 /= "111111110001011101111110001" OR uut_h_1_1 /= "111111111010100010101000011" OR uut_h_1_2 /= "111111110101011000101111100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0000000";
              state <= "1100111";
            ELSE
              state <= "0000100";
            END IF;
            uut_rst <= '0';
          WHEN "0000100" =>
            uut_h_0_0_i <= "111111110001111100010100101";
            uut_h_0_1_i <= "000000000111011111100110011";
            uut_h_0_2_i <= "000000001001000011000001110";
            uut_h_1_0_i <= "111111111100011110010111011";
            uut_h_1_1_i <= "111111110011010101011010111";
            uut_h_1_2_i <= "000000000001000010010110011";
            uut_xb <= "111111110010010001010100001";
            uut_yb <= "000000000100000001101001010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000110111010111111110" OR uut_h_0_1 /= "000000001111011110000010111" OR uut_h_0_2 /= "111111111110000100111010111" OR uut_h_1_0 /= "000000001101011110111001011" OR uut_h_1_1 /= "000000001100101011101000101" OR uut_h_1_2 /= "000000001100110101110010000" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0000001";
              state <= "1100111";
            ELSE
              state <= "0000101";
            END IF;
            uut_rst <= '0';
          WHEN "0000101" =>
            uut_h_0_0_i <= "111111110000110010100011000";
            uut_h_0_1_i <= "111111111110011010110110111";
            uut_h_0_2_i <= "111111111111111100110100001";
            uut_h_1_0_i <= "111111110001111111000100000";
            uut_h_1_1_i <= "000000000101100000111100011";
            uut_h_1_2_i <= "111111110001100011111010010";
            uut_xb <= "000000000100100010000011111";
            uut_yb <= "000000001001001010100001010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001011101001011001100" OR uut_h_0_1 /= "111111110010010000111010000" OR uut_h_0_2 /= "111111111000110110101010110" OR uut_h_1_0 /= "111111111000110010011000001" OR uut_h_1_1 /= "111111111100000111110001000" OR uut_h_1_2 /= "000000001010110000110010010" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0000010";
              state <= "1100111";
            ELSE
              state <= "0000110";
            END IF;
            uut_rst <= '0';
          WHEN "0000110" =>
            uut_h_0_0_i <= "111111111001010000001011100";
            uut_h_0_1_i <= "000000000011000010110100101";
            uut_h_0_2_i <= "111111111101001011001001000";
            uut_h_1_0_i <= "111111111111111011101000100";
            uut_h_1_1_i <= "000000000001001010100110001";
            uut_h_1_2_i <= "000000001001011010000111111";
            uut_xb <= "111111111110110011011010110";
            uut_yb <= "111111111011110001010011011";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000111101000101010111" OR uut_h_0_1 /= "000000000010011100100100101" OR uut_h_0_2 /= "000000000101100010010110100" OR uut_h_1_0 /= "111111110000011010000111111" OR uut_h_1_1 /= "000000001001110101100000110" OR uut_h_1_2 /= "000000000110111000000110010" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0000011";
              state <= "1100111";
            ELSE
              state <= "0000111";
            END IF;
            uut_rst <= '0';
          WHEN "0000111" =>
            uut_h_0_0_i <= "000000000101101111110000101";
            uut_h_0_1_i <= "111111111111101101110011010";
            uut_h_0_2_i <= "111111110010001000010111110";
            uut_h_1_0_i <= "000000000010001010110011111";
            uut_h_1_1_i <= "111111111100110000000010101";
            uut_h_1_2_i <= "111111111101001001110010010";
            uut_xb <= "000000001000111110111010101";
            uut_yb <= "000000000111010101000001110";
            uut_input_valid <= '0';
            IF uut_h_0_0 /= "111111110001111100010100101" OR uut_h_0_1 /= "000000000111011111100110011" OR uut_h_0_2 /= "111111101101010111101010110" OR uut_h_1_0 /= "111111111100011110010111011" OR uut_h_1_1 /= "111111110011010101011010111" OR uut_h_1_2 /= "000000000101001110010100111" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0000100";
              state <= "1100111";
            ELSE
              state <= "0001000";
            END IF;
            uut_rst <= '0';
          WHEN "0001000" =>
            uut_h_0_0_i <= "000000001000100000000011010";
            uut_h_0_1_i <= "000000001000101001010001111";
            uut_h_0_2_i <= "111111111100101011001010100";
            uut_h_1_0_i <= "000000001000001101011110100";
            uut_h_1_1_i <= "000000001111010100010011000";
            uut_h_1_2_i <= "111111111111101111101111010";
            uut_xb <= "111111110001001011101101001";
            uut_yb <= "000000001111001011100010000";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110000110010100011000" OR uut_h_0_1 /= "111111111110011010110110111" OR uut_h_0_2 /= "000000001001101100100011011" OR uut_h_1_0 /= "111111110001111111000100000" OR uut_h_1_1 /= "000000000101100000111100011" OR uut_h_1_2 /= "111111111011100010010110000" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0000101";
              state <= "1100111";
            ELSE
              state <= "0001001";
            END IF;
            uut_rst <= '0';
          WHEN "0001001" =>
            uut_h_0_0_i <= "000000000111001111101110000";
            uut_h_0_1_i <= "000000000110100011011110101";
            uut_h_0_2_i <= "111111111101001001011001101";
            uut_h_1_0_i <= "111111110100101111000010000";
            uut_h_1_1_i <= "111111111100001100010001100";
            uut_h_1_2_i <= "111111110100100100110110000";
            uut_xb <= "000000001101110001001001011";
            uut_yb <= "111111110000001001101010100";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111001010000001011100" OR uut_h_0_1 /= "000000000011000010110100101" OR uut_h_0_2 /= "111111111100010001110001001" OR uut_h_1_0 /= "111111111111111011101000100" OR uut_h_1_1 /= "000000000001001010100110001" OR uut_h_1_2 /= "000000000101011110110100100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0000110";
              state <= "1100111";
            ELSE
              state <= "0001010";
            END IF;
            uut_rst <= '0';
          WHEN "0001010" =>
            uut_h_0_0_i <= "000000000100110011010010000";
            uut_h_0_1_i <= "000000001010111110110101011";
            uut_h_0_2_i <= "111111110010111111000101111";
            uut_h_1_0_i <= "000000000101101101101000100";
            uut_h_1_1_i <= "111111111001011010000001110";
            uut_h_1_2_i <= "000000001001100010000100011";
            uut_xb <= "000000001001000100011010101";
            uut_yb <= "000000000011111101110010110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000101101111110000101" OR uut_h_0_1 /= "111111111111101101110011010" OR uut_h_0_2 /= "111111111000000001001001100" OR uut_h_1_0 /= "000000000010001010110011111" OR uut_h_1_1 /= "111111111100110000000010101" OR uut_h_1_2 /= "000000000100110000001000100" OR uut_output_valid /= '0' THEN
              FAIL <= '1';
              FAIL_NUM <= "0000111";
              state <= "1100111";
            ELSE
              state <= "0001011";
            END IF;
            uut_rst <= '0';
          WHEN "0001011" =>
            uut_h_0_0_i <= "000000001010011010011100110";
            uut_h_0_1_i <= "111111110111111111010100100";
            uut_h_0_2_i <= "111111111000111110110101111";
            uut_h_1_0_i <= "111111110001000111101110011";
            uut_h_1_1_i <= "111111111111011000111000000";
            uut_h_1_2_i <= "000000000011001011000010110";
            uut_xb <= "111111110100111101110110001";
            uut_yb <= "000000001010101011110110010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001000100000000011010" OR uut_h_0_1 /= "000000001000101001010001111" OR uut_h_0_2 /= "111111101101100001110001010" OR uut_h_1_0 /= "000000001000001101011110100" OR uut_h_1_1 /= "000000001111010100010011000" OR uut_h_1_2 /= "000000000111111111110101010" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0001000";
              state <= "1100111";
            ELSE
              state <= "0001100";
            END IF;
            uut_rst <= '0';
          WHEN "0001100" =>
            uut_h_0_0_i <= "111111110110001111001001000";
            uut_h_0_1_i <= "000000000101011110011100100";
            uut_h_0_2_i <= "111111111111111110111100000";
            uut_h_1_0_i <= "000000001010100011011001111";
            uut_h_1_1_i <= "111111110001101011001111110";
            uut_h_1_2_i <= "000000001110001011111000001";
            uut_xb <= "111111111100000011001100100";
            uut_yb <= "111111110011101000111110001";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000111001111101110000" OR uut_h_0_1 /= "000000000110100011011110101" OR uut_h_0_2 /= "000000001011001011000010101" OR uut_h_1_0 /= "111111110100101111000010000" OR uut_h_1_1 /= "111111111100001100010001100" OR uut_h_1_2 /= "111111101010101001011110010" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0001001";
              state <= "1100111";
            ELSE
              state <= "0001101";
            END IF;
            uut_rst <= '0';
          WHEN "0001101" =>
            uut_h_0_0_i <= "000000001110111000000000111";
            uut_h_0_1_i <= "000000000110111011110000001";
            uut_h_0_2_i <= "000000001000000111001101111";
            uut_h_1_0_i <= "111111111101110101110010001";
            uut_h_1_1_i <= "000000000000001101111001101";
            uut_h_1_2_i <= "000000001010110000001000111";
            uut_xb <= "000000000001000110100000001";
            uut_yb <= "111111111101111011001101111";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000100110011010010000" OR uut_h_0_1 /= "000000001010111110110101011" OR uut_h_0_2 /= "111111110110100111001001010" OR uut_h_1_0 /= "000000000101101101101000100" OR uut_h_1_1 /= "111111111001011010000001110" OR uut_h_1_2 /= "000000001011111001001100111" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0001010";
              state <= "1100111";
            ELSE
              state <= "0001110";
            END IF;
            uut_rst <= '0';
          WHEN "0001110" =>
            uut_h_0_0_i <= "111111110101000010111110100";
            uut_h_0_1_i <= "111111110011011100101100001";
            uut_h_0_2_i <= "111111111101101011001110011";
            uut_h_1_0_i <= "000000000011001101110010010";
            uut_h_1_1_i <= "000000001100110011001010010";
            uut_h_1_2_i <= "111111110100111000000100110";
            uut_xb <= "111111111110010100001101100";
            uut_yb <= "000000000001000011001000111";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001010011010011100110" OR uut_h_0_1 /= "111111110111111111010100100" OR uut_h_0_2 /= "111111111010011110101001110" OR uut_h_1_0 /= "111111110001000111101110011" OR uut_h_1_1 /= "111111111111011000111000000" OR uut_h_1_2 /= "000000000100000000010101000" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0001011";
              state <= "1100111";
            ELSE
              state <= "0001111";
            END IF;
            uut_rst <= '0';
          WHEN "0001111" =>
            uut_h_0_0_i <= "111111111011010110010100110";
            uut_h_0_1_i <= "000000000111011111011010111";
            uut_h_0_2_i <= "000000000100100000111110111";
            uut_h_1_0_i <= "000000001000101111010101101";
            uut_h_1_1_i <= "111111111101000000010111111";
            uut_h_1_2_i <= "111111110100000101000011010";
            uut_xb <= "111111111001111011110101110";
            uut_yb <= "000000000010100000111010111";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110110001111001001000" OR uut_h_0_1 /= "000000000101011110011100100" OR uut_h_0_2 /= "111111111101110110100101100" OR uut_h_1_0 /= "000000001010100011011001111" OR uut_h_1_1 /= "111111110001101011001111110" OR uut_h_1_2 /= "111111111001010111011010010" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0001100";
              state <= "1100111";
            ELSE
              state <= "0010000";
            END IF;
            uut_rst <= '0';
          WHEN "0010000" =>
            uut_h_0_0_i <= "000000001110001100100000101";
            uut_h_0_1_i <= "000000001101101111011110110";
            uut_h_0_2_i <= "111111111000010100011101010";
            uut_h_1_0_i <= "111111111101101010010111110";
            uut_h_1_1_i <= "000000001101100110010111010";
            uut_h_1_2_i <= "000000001001001011011111010";
            uut_xb <= "000000000010000000000011100";
            uut_yb <= "000000000101111010011101010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001110111000000000111" OR uut_h_0_1 /= "000000000110111011110000001" OR uut_h_0_2 /= "000000001001000101101101111" OR uut_h_1_0 /= "111111111101110101110010001" OR uut_h_1_1 /= "000000000000001101111001101" OR uut_h_1_2 /= "000000001000110110101011010" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0001101";
              state <= "1100111";
            ELSE
              state <= "0010001";
            END IF;
            uut_rst <= '0';
          WHEN "0010001" =>
            uut_h_0_0_i <= "111111110010111101001110100";
            uut_h_0_1_i <= "111111110011000101110100110";
            uut_h_0_2_i <= "111111110000010111001110100";
            uut_h_1_0_i <= "000000001011111011000010101";
            uut_h_1_1_i <= "000000001011000100010111100";
            uut_h_1_2_i <= "000000000000110000100000001";
            uut_xb <= "111111111100010100110001110";
            uut_yb <= "000000000100110001110001010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110101000010111110100" OR uut_h_0_1 /= "111111110011011100101100001" OR uut_h_0_2 /= "111111111011101010010100001" OR uut_h_1_0 /= "000000000011001101110010010" OR uut_h_1_1 /= "000000001100110011001010010" OR uut_h_1_2 /= "111111110101011011001010110" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0001110";
              state <= "1100111";
            ELSE
              state <= "0010010";
            END IF;
            uut_rst <= '0';
          WHEN "0010010" =>
            uut_h_0_0_i <= "000000001000011010010100101";
            uut_h_0_1_i <= "111111111000111001110000110";
            uut_h_0_2_i <= "000000000100001101100100000";
            uut_h_1_0_i <= "000000000010011011000000010";
            uut_h_1_1_i <= "000000001010110111111111000";
            uut_h_1_2_i <= "000000001010101010111100001";
            uut_xb <= "111111111100110100110101110";
            uut_yb <= "000000000001101111000111010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111011010110010100110" OR uut_h_0_1 /= "000000000111011111011010111" OR uut_h_0_2 /= "111111111011100000101001011" OR uut_h_1_0 /= "000000001000101111010101101" OR uut_h_1_1 /= "111111111101000000010111111" OR uut_h_1_2 /= "111111111010011000000111001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0001111";
              state <= "1100111";
            ELSE
              state <= "0010011";
            END IF;
            uut_rst <= '0';
          WHEN "0010011" =>
            uut_h_0_0_i <= "111111111110001101000010010";
            uut_h_0_1_i <= "111111110001000010110010111";
            uut_h_0_2_i <= "000000001111001110011011110";
            uut_h_1_0_i <= "111111110010111001000110110";
            uut_h_1_1_i <= "111111111101110000000111001";
            uut_h_1_2_i <= "000000000000101101110000001";
            uut_xb <= "111111111100010000111001000";
            uut_yb <= "000000001100010011010110111";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001110001100100000101" OR uut_h_0_1 /= "000000001101101111011110110" OR uut_h_0_2 /= "111111110011011101110110111" OR uut_h_1_0 /= "111111111101101010010111110" OR uut_h_1_1 /= "000000001101100110010111010" OR uut_h_1_2 /= "000000001010010110111111000" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0010000";
              state <= "1100111";
            ELSE
              state <= "0010100";
            END IF;
            uut_rst <= '0';
          WHEN "0010100" =>
            uut_h_0_0_i <= "111111111000001010010001101";
            uut_h_0_1_i <= "111111111100110000001010011";
            uut_h_0_2_i <= "000000001100100111111101011";
            uut_h_1_0_i <= "000000001101000101101110111";
            uut_h_1_1_i <= "000000000100000000000010100";
            uut_h_1_2_i <= "111111110110110110100111001";
            uut_xb <= "000000001100001011011011100";
            uut_yb <= "111111110111100001100001110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110010111101001110100" OR uut_h_0_1 /= "111111110011000101110100110" OR uut_h_0_2 /= "111111101101100010111100110" OR uut_h_1_0 /= "000000001011111011000010101" OR uut_h_1_1 /= "000000001011000100010111100" OR uut_h_1_2 /= "000000000100111110000010000" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0010001";
              state <= "1100111";
            ELSE
              state <= "0010101";
            END IF;
            uut_rst <= '0';
          WHEN "0010101" =>
            uut_h_0_0_i <= "111111110111110101011110111";
            uut_h_0_1_i <= "000000001010011010110111110";
            uut_h_0_2_i <= "111111111100100000010110010";
            uut_h_1_0_i <= "000000000100100000100110010";
            uut_h_1_1_i <= "000000001100010001110010110";
            uut_h_1_2_i <= "000000001001101001000110100";
            uut_xb <= "000000000100000000010101101";
            uut_yb <= "000000000110010111100001011";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001000011010010100101" OR uut_h_0_1 /= "111111111000111001110000110" OR uut_h_0_2 /= "000000000011011110011111101" OR uut_h_1_0 /= "000000000010011011000000010" OR uut_h_1_1 /= "000000001010110111111111000" OR uut_h_1_2 /= "000000001011101101010010011" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0010010";
              state <= "1100111";
            ELSE
              state <= "0010110";
            END IF;
            uut_rst <= '0';
          WHEN "0010110" =>
            uut_h_0_0_i <= "111111110010101111110111000";
            uut_h_0_1_i <= "111111111000011011111111001";
            uut_h_0_2_i <= "111111111111110110110111011";
            uut_h_1_0_i <= "000000000000111111110110110";
            uut_h_1_1_i <= "111111110111100000110101110";
            uut_h_1_2_i <= "111111110100111000000010111";
            uut_xb <= "000000000101000011011111010";
            uut_yb <= "000000000010000000111010110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111110001101000010010" OR uut_h_0_1 /= "111111110001000010110010111" OR uut_h_0_2 /= "000000010110100100011110110" OR uut_h_1_0 /= "111111110010111001000110110" OR uut_h_1_1 /= "111111111101110000000111001" OR uut_h_1_2 /= "000000001011101011110111001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0010011";
              state <= "1100111";
            ELSE
              state <= "0010111";
            END IF;
            uut_rst <= '0';
          WHEN "0010111" =>
            uut_h_0_0_i <= "111111111001010101101010100";
            uut_h_0_1_i <= "111111111000111110111011111";
            uut_h_0_2_i <= "000000001001000000010010100";
            uut_h_1_0_i <= "000000000011111010011110110";
            uut_h_1_1_i <= "111111111101001100010101011";
            uut_h_1_2_i <= "111111110100010101011110100";
            uut_xb <= "111111111001010001001011001";
            uut_yb <= "111111111111111111000110000";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111000001010010001101" OR uut_h_0_1 /= "111111111100110000001010011" OR uut_h_0_2 /= "000000011101000011001011100" OR uut_h_1_0 /= "000000001101000101101110111" OR uut_h_1_1 /= "000000000100000000000010100" OR uut_h_1_2 /= "111111100110100010001000011" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0010100";
              state <= "1100111";
            ELSE
              state <= "0011000";
            END IF;
            uut_rst <= '0';
          WHEN "0011000" =>
            uut_h_0_0_i <= "000000001001000100110010110";
            uut_h_0_1_i <= "000000000110010010101011010";
            uut_h_0_2_i <= "000000001100010111010111110";
            uut_h_1_0_i <= "000000000101101010100111111";
            uut_h_1_1_i <= "111111110100001000001101111";
            uut_h_1_2_i <= "000000000000011110101110101";
            uut_xb <= "000000001111010000011110010";
            uut_yb <= "111111110100000000111100010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110111110101011110111" OR uut_h_0_1 /= "000000001010011010110111110" OR uut_h_0_2 /= "111111111110011010000110000" OR uut_h_1_0 /= "000000000100100000100110010" OR uut_h_1_1 /= "000000001100010001110010110" OR uut_h_1_2 /= "000000001001111111101010001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0010101";
              state <= "1100111";
            ELSE
              state <= "0011001";
            END IF;
            uut_rst <= '0';
          WHEN "0011001" =>
            uut_h_0_0_i <= "000000001000000100100110000";
            uut_h_0_1_i <= "111111110110000110111011010";
            uut_h_0_2_i <= "111111111010011010001011110";
            uut_h_1_0_i <= "000000001010011101110011010";
            uut_h_1_1_i <= "111111111101101101110110111";
            uut_h_1_2_i <= "111111110100010011110111101";
            uut_xb <= "000000000010010100000001001";
            uut_yb <= "000000001001010110000100000";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110010101111110111000" OR uut_h_0_1 /= "111111111000011011111111001" OR uut_h_0_2 /= "000000001010000011001110011" OR uut_h_1_0 /= "000000000000111111110110110" OR uut_h_1_1 /= "111111110111100000110101110" OR uut_h_1_2 /= "111111110111101001001011001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0010110";
              state <= "1100111";
            ELSE
              state <= "0011010";
            END IF;
            uut_rst <= '0';
          WHEN "0011010" =>
            uut_h_0_0_i <= "111111111101011011100111101";
            uut_h_0_1_i <= "000000001100110001010100011";
            uut_h_0_2_i <= "111111110001101010001001000";
            uut_h_1_0_i <= "000000000001000010101000101";
            uut_h_1_1_i <= "000000000001011011110100011";
            uut_h_1_2_i <= "000000001001111000000001001";
            uut_xb <= "111111110111010100010101111";
            uut_yb <= "000000001010010100010001110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111001010101101010100" OR uut_h_0_1 /= "111111111000111110111011111" OR uut_h_0_2 /= "111111111111011101101100100" OR uut_h_1_0 /= "000000000011111010011110110" OR uut_h_1_1 /= "111111111101001100010101011" OR uut_h_1_2 /= "111111110101111101110011000" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0010111";
              state <= "1100111";
            ELSE
              state <= "0011011";
            END IF;
            uut_rst <= '0';
          WHEN "0011011" =>
            uut_h_0_0_i <= "111111111011001001001011110";
            uut_h_0_1_i <= "000000001110100100100110001";
            uut_h_0_2_i <= "000000001110000011010000110";
            uut_h_1_0_i <= "111111110101010010111000100";
            uut_h_1_1_i <= "000000000101110001001111000";
            uut_h_1_2_i <= "000000000101110001000010011";
            uut_xb <= "111111111000001101101101000";
            uut_yb <= "000000001100010101101111101";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001001000100110010110" OR uut_h_0_1 /= "000000000110010010101011010" OR uut_h_0_2 /= "000000010111101011101001010" OR uut_h_1_0 /= "000000000101101010100111111" OR uut_h_1_1 /= "111111110100001000001101111" OR uut_h_1_2 /= "111111100110001100101111011" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0011000";
              state <= "1100111";
            ELSE
              state <= "0011100";
            END IF;
            uut_rst <= '0';
          WHEN "0011100" =>
            uut_h_0_0_i <= "000000001101011100001111110";
            uut_h_0_1_i <= "000000001000100011101000011";
            uut_h_0_2_i <= "111111111110010101010001110";
            uut_h_1_0_i <= "111111111001100110100001111";
            uut_h_1_1_i <= "111111110010101101111110110";
            uut_h_1_2_i <= "000000000100110101110000011";
            uut_xb <= "000000000001000000011010000";
            uut_yb <= "000000000100010010000001100";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001000000100100110000" OR uut_h_0_1 /= "111111110110000110111011010" OR uut_h_0_2 /= "000000000001010101010001100" OR uut_h_1_0 /= "000000001010011101110011010" OR uut_h_1_1 /= "111111111101101101110110111" OR uut_h_1_2 /= "111111111101011110011110000" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0011001";
              state <= "1100111";
            ELSE
              state <= "0011101";
            END IF;
            uut_rst <= '0';
          WHEN "0011101" =>
            uut_h_0_0_i <= "111111110000011100110111100";
            uut_h_0_1_i <= "111111110011101001100001111";
            uut_h_0_2_i <= "111111111001011011101100011";
            uut_h_1_0_i <= "111111111111000011010100100";
            uut_h_1_1_i <= "111111111110001010010100110";
            uut_h_1_2_i <= "000000001110011010010110101";
            uut_xb <= "111111110110100111100010100";
            uut_yb <= "000000000001110000001001110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111101011011100111101" OR uut_h_0_1 /= "000000001100110001010100011" OR uut_h_0_2 /= "111111011111010110010001110" OR uut_h_1_0 /= "000000000001000010101000101" OR uut_h_1_1 /= "000000000001011011110100011" OR uut_h_1_2 /= "000000010011110101010000001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0011010";
              state <= "1100111";
            ELSE
              state <= "0011110";
            END IF;
            uut_rst <= '0';
          WHEN "0011110" =>
            uut_h_0_0_i <= "000000001100001000110000110";
            uut_h_0_1_i <= "000000001100101000110000011";
            uut_h_0_2_i <= "111111110110000011011000110";
            uut_h_1_0_i <= "000000000001110110011111100";
            uut_h_1_1_i <= "000000001010111100000110001";
            uut_h_1_2_i <= "111111110100111010101001111";
            uut_xb <= "111111110000010010100110110";
            uut_yb <= "000000000011000101100010000";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111011001001001011110" OR uut_h_0_1 /= "000000001110100100100110001" OR uut_h_0_2 /= "111111111000101010011110000" OR uut_h_1_0 /= "111111110101010010111000100" OR uut_h_1_1 /= "000000000101110001001111000" OR uut_h_1_2 /= "000000001000011100101000001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0011011";
              state <= "1100111";
            ELSE
              state <= "0011111";
            END IF;
            uut_rst <= '0';
          WHEN "0011111" =>
            uut_h_0_0_i <= "000000000011011111010101010";
            uut_h_0_1_i <= "111111111001101000101111111";
            uut_h_0_2_i <= "000000000111011100111000101";
            uut_h_1_0_i <= "000000001101011001111101001";
            uut_h_1_1_i <= "111111111111110110111011111";
            uut_h_1_2_i <= "111111110011101111001000000";
            uut_xb <= "000000001001111010011100101";
            uut_yb <= "000000000111110110001111010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001101011100001111110" OR uut_h_0_1 /= "000000001000100011101000011" OR uut_h_0_2 /= "111111111100001101000010001" OR uut_h_1_0 /= "111111111001100110100001111" OR uut_h_1_1 /= "111111110010101101111110110" OR uut_h_1_2 /= "000000001101000101000000001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0011100";
              state <= "1100111";
            ELSE
              state <= "0100000";
            END IF;
            uut_rst <= '0';
          WHEN "0100000" =>
            uut_h_0_0_i <= "111111111010110010011110000";
            uut_h_0_1_i <= "111111110010110010101110000";
            uut_h_0_2_i <= "111111111000100011011110110";
            uut_h_1_0_i <= "000000000010101100101100101";
            uut_h_1_1_i <= "000000001010100001001101101";
            uut_h_1_2_i <= "000000001111000001100000001";
            uut_xb <= "111111111001100110010001110";
            uut_yb <= "111111111101001010000110110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110000011100110111100" OR uut_h_0_1 /= "111111110011101001100001111" OR uut_h_0_2 /= "111111101000010010010001101" OR uut_h_1_0 /= "111111111111000011010100100" OR uut_h_1_1 /= "111111111110001010010100110" OR uut_h_1_2 /= "000000001111110011110100001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0011101";
              state <= "1100111";
            ELSE
              state <= "0100001";
            END IF;
            uut_rst <= '0';
          WHEN "0100001" =>
            uut_h_0_0_i <= "111111110111100100010101000";
            uut_h_0_1_i <= "111111110101110001110000110";
            uut_h_0_2_i <= "111111111110110011110001101";
            uut_h_1_0_i <= "111111110110001111011110010";
            uut_h_1_1_i <= "000000000000101101101111001";
            uut_h_1_2_i <= "000000001101100110111000000";
            uut_xb <= "111111110000000010000100001";
            uut_yb <= "000000001101000000101110101";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001100001000110000110" OR uut_h_0_1 /= "000000001100101000110000011" OR uut_h_0_2 /= "111111101111110100101000011" OR uut_h_1_0 /= "000000000001110110011111100" OR uut_h_1_1 /= "000000001010111100000110001" OR uut_h_1_2 /= "111111110111101101011110100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0011110";
              state <= "1100111";
            ELSE
              state <= "0100010";
            END IF;
            uut_rst <= '0';
          WHEN "0100010" =>
            uut_h_0_0_i <= "000000000101110000101110011";
            uut_h_0_1_i <= "111111110011010010110001101";
            uut_h_0_2_i <= "000000000100000000011111110";
            uut_h_1_0_i <= "000000000000011110100111110";
            uut_h_1_1_i <= "000000001111111001100111000";
            uut_h_1_2_i <= "111111111100100101100111010";
            uut_xb <= "000000000001011100101111100";
            uut_yb <= "000000000000010010101010000";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000011011111010101010" OR uut_h_0_1 /= "111111111001101000101111111" OR uut_h_0_2 /= "000000010010010100101101001" OR uut_h_1_0 /= "000000001101011001111101001" OR uut_h_1_1 /= "111111111111110110111011111" OR uut_h_1_2 /= "111111110011010110001111100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0011111";
              state <= "1100111";
            ELSE
              state <= "0100011";
            END IF;
            uut_rst <= '0';
          WHEN "0100011" =>
            uut_h_0_0_i <= "111111110111111001011001110";
            uut_h_0_1_i <= "111111110001100010110100001";
            uut_h_0_2_i <= "000000001111000111011110011";
            uut_h_1_0_i <= "111111110001011100111110000";
            uut_h_1_1_i <= "111111111010000111110100110";
            uut_h_1_2_i <= "000000000010110001000101000";
            uut_xb <= "000000000111010010010100110";
            uut_yb <= "000000000100110101001110001";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111010110010011110000" OR uut_h_0_1 /= "111111110010110010101110000" OR uut_h_0_2 /= "111111101101101110001010001" OR uut_h_1_0 /= "000000000010101100101100101" OR uut_h_1_1 /= "000000001010100001001101101" OR uut_h_1_2 /= "000000001111001000010010101" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0100000";
              state <= "1100111";
            ELSE
              state <= "0100100";
            END IF;
            uut_rst <= '0';
          WHEN "0100100" =>
            uut_h_0_0_i <= "000000000101010001001000011";
            uut_h_0_1_i <= "111111111100110000000000010";
            uut_h_0_2_i <= "111111110100010000001000000";
            uut_h_1_0_i <= "000000001110000010100111101";
            uut_h_1_1_i <= "000000000101011101000110001";
            uut_h_1_2_i <= "111111111110000011011111010";
            uut_xb <= "111111111100101001001111010";
            uut_yb <= "111111111100101111101010010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110111100100010101000" OR uut_h_0_1 /= "111111110101110001110000110" OR uut_h_0_2 /= "111111101110101111010010110" OR uut_h_1_0 /= "111111110110001111011110010" OR uut_h_1_1 /= "000000000000101101101111001" OR uut_h_1_2 /= "000000010000010011001001010" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0100001";
              state <= "1100111";
            ELSE
              state <= "0100101";
            END IF;
            uut_rst <= '0';
          WHEN "0100101" =>
            uut_h_0_0_i <= "000000001000000010110000110";
            uut_h_0_1_i <= "111111110010110101100111010";
            uut_h_0_2_i <= "000000000100011010100010110";
            uut_h_1_0_i <= "000000000000101101110001100";
            uut_h_1_1_i <= "111111111000000001101111101";
            uut_h_1_2_i <= "000000000110101100111100011";
            uut_xb <= "000000001101110101001000101";
            uut_yb <= "111111110010111100111000101";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000101110000101110011" OR uut_h_0_1 /= "111111110011010010110001101" OR uut_h_0_2 /= "000000000101001010101010010" OR uut_h_1_0 /= "000000000000011110100111110" OR uut_h_1_1 /= "000000001111111001100111000" OR uut_h_1_2 /= "111111111100100010111101011" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0100010";
              state <= "1100111";
            ELSE
              state <= "0100110";
            END IF;
            uut_rst <= '0';
          WHEN "0100110" =>
            uut_h_0_0_i <= "000000001110100000110110011";
            uut_h_0_1_i <= "000000000011000110101010110";
            uut_h_0_2_i <= "111111111001100110011111000";
            uut_h_1_0_i <= "111111110101001101011001111";
            uut_h_1_1_i <= "111111110111101011111111000";
            uut_h_1_2_i <= "000000001010000010001000111";
            uut_xb <= "111111111011010101111101011";
            uut_yb <= "111111110100001110010110111";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110111111001011001110" OR uut_h_0_1 /= "111111110001100010110100001" OR uut_h_0_2 /= "000000011110011101010110011" OR uut_h_1_0 /= "111111110001011100111110000" OR uut_h_1_1 /= "111111111010000111110100110" OR uut_h_1_2 /= "000000001111111111111000100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0100011";
              state <= "1100111";
            ELSE
              state <= "0100111";
            END IF;
            uut_rst <= '0';
          WHEN "0100111" =>
            uut_h_0_0_i <= "111111110101000011111100111";
            uut_h_0_1_i <= "111111110010110001000111010";
            uut_h_0_2_i <= "000000000100110110000100011";
            uut_h_1_0_i <= "111111110001111111010001101";
            uut_h_1_1_i <= "000000000011101111001011100";
            uut_h_1_2_i <= "111111111111111101010101001";
            uut_xb <= "000000001010100100111111001";
            uut_yb <= "000000001010001100000000000";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000101010001001000011" OR uut_h_0_1 /= "111111111100110000000000010" OR uut_h_0_2 /= "111111110001010101110000010" OR uut_h_1_0 /= "000000001110000010100111101" OR uut_h_1_1 /= "000000000101011101000110001" OR uut_h_1_2 /= "111111111110110110101001001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0100100";
              state <= "1100111";
            ELSE
              state <= "0101000";
            END IF;
            uut_rst <= '0';
          WHEN "0101000" =>
            uut_h_0_0_i <= "000000001110000001010111101";
            uut_h_0_1_i <= "111111110000001111000100001";
            uut_h_0_2_i <= "111111111011101111110101101";
            uut_h_1_0_i <= "111111110000000000101010101";
            uut_h_1_1_i <= "111111110011011001111100110";
            uut_h_1_2_i <= "111111110111101010101101110";
            uut_xb <= "111111110111111111001110001";
            uut_yb <= "111111111100011000101101010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001000000010110000110" OR uut_h_0_1 /= "111111110010110101100111010" OR uut_h_0_2 /= "000000000000100011101110011" OR uut_h_1_0 /= "000000000000101101110001100" OR uut_h_1_1 /= "111111111000000001101111101" OR uut_h_1_2 /= "111111110010100010001000010" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0100101";
              state <= "1100111";
            ELSE
              state <= "0101001";
            END IF;
            uut_rst <= '0';
          WHEN "0101001" =>
            uut_h_0_0_i <= "111111111101011110010010010";
            uut_h_0_1_i <= "111111111000101000111100101";
            uut_h_0_2_i <= "000000001010011011110110110";
            uut_h_1_0_i <= "000000000100011110111000001";
            uut_h_1_1_i <= "000000001011000000011110011";
            uut_h_1_2_i <= "111111110101110101001000010";
            uut_xb <= "000000000011100001111111110";
            uut_yb <= "000000000110011100110001111";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001110100000110110011" OR uut_h_0_1 /= "000000000011000110101010110" OR uut_h_0_2 /= "111111111011011101000000100" OR uut_h_1_0 /= "111111110101001101011001111" OR uut_h_1_1 /= "111111110111101011111111000" OR uut_h_1_2 /= "111111110100111111111100100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0100110";
              state <= "1100111";
            ELSE
              state <= "0101010";
            END IF;
            uut_rst <= '0';
          WHEN "0101010" =>
            uut_h_0_0_i <= "111111110011100100100101111";
            uut_h_0_1_i <= "000000001001111111011100111";
            uut_h_0_2_i <= "000000000111011001101010001";
            uut_h_1_0_i <= "111111110011000100001111110";
            uut_h_1_1_i <= "000000001010000100010000011";
            uut_h_1_2_i <= "000000001100111011000110010";
            uut_xb <= "111111110010010000110001001";
            uut_yb <= "111111110111101110001000110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110101000011111100111" OR uut_h_0_1 /= "111111110010110001000111010" OR uut_h_0_2 /= "000000011111000101000110100" OR uut_h_1_0 /= "111111110001111111010001101" OR uut_h_1_1 /= "000000000011101111001011100" OR uut_h_1_2 /= "000000010001000001111000101" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0100111";
              state <= "1100111";
            ELSE
              state <= "0101011";
            END IF;
            uut_rst <= '0';
          WHEN "0101011" =>
            uut_h_0_0_i <= "000000000111011010110111000";
            uut_h_0_1_i <= "000000000001010010010111000";
            uut_h_0_2_i <= "111111110011101110001111111";
            uut_h_1_0_i <= "111111110001010010111011010";
            uut_h_1_1_i <= "000000001110100001011100000";
            uut_h_1_2_i <= "000000000100101011011101010";
            uut_xb <= "000000001111011110001100111";
            uut_yb <= "111111110111111100100110111";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001110000001010111101" OR uut_h_0_1 /= "111111110000001111000100001" OR uut_h_0_2 /= "111111110111001100100010100" OR uut_h_1_0 /= "111111110000000000101010101" OR uut_h_1_1 /= "111111110011011001111100110" OR uut_h_1_2 /= "111111101001001100111010100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0101000";
              state <= "1100111";
            ELSE
              state <= "0101100";
            END IF;
            uut_rst <= '0';
          WHEN "0101100" =>
            uut_h_0_0_i <= "000000000011011001110100010";
            uut_h_0_1_i <= "111111111111101001100011010";
            uut_h_0_2_i <= "000000001100110101001100100";
            uut_h_1_0_i <= "000000001010001000100101111";
            uut_h_1_1_i <= "000000001000010101111110001";
            uut_h_1_2_i <= "111111110110110110110000100";
            uut_xb <= "000000001001000111000101011";
            uut_yb <= "111111110110001110001101110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111101011110010010010" OR uut_h_0_1 /= "111111111000101000111100101" OR uut_h_0_2 /= "000000010001011111011011011" OR uut_h_1_0 /= "000000000100011110111000001" OR uut_h_1_1 /= "000000001011000000011110011" OR uut_h_1_2 /= "111111110110110110100111101" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0101001";
              state <= "1100111";
            ELSE
              state <= "0101101";
            END IF;
            uut_rst <= '0';
          WHEN "0101101" =>
            uut_h_0_0_i <= "000000000111111001101000010";
            uut_h_0_1_i <= "111111111000010101100110100";
            uut_h_0_2_i <= "000000001101010110010001111";
            uut_h_1_0_i <= "111111111111001101111100010";
            uut_h_1_1_i <= "111111110010101101101101110";
            uut_h_1_2_i <= "111111111111000011100111110";
            uut_xb <= "000000001000011010100100000";
            uut_yb <= "000000001000101101011010001";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110011100100100101111" OR uut_h_0_1 /= "000000001001111111011100111" OR uut_h_0_2 /= "111111110100001010010110011" OR uut_h_1_0 /= "111111110011000100001111110" OR uut_h_1_1 /= "000000001010000100010000011" OR uut_h_1_2 /= "111111111110101111110111110" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0101010";
              state <= "1100111";
            ELSE
              state <= "0101110";
            END IF;
            uut_rst <= '0';
          WHEN "0101110" =>
            uut_h_0_0_i <= "111111110000101011100111110";
            uut_h_0_1_i <= "111111111010010111111000111";
            uut_h_0_2_i <= "000000001101110000100010101";
            uut_h_1_0_i <= "000000001100001010001101100";
            uut_h_1_1_i <= "000000000101011010001100111";
            uut_h_1_2_i <= "111111111001000001011101000";
            uut_xb <= "000000000111110110000110011";
            uut_yb <= "111111111111010001001010111";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000111011010110111000" OR uut_h_0_1 /= "000000000001010010010111000" OR uut_h_0_2 /= "111111111100101010101101111" OR uut_h_1_0 /= "111111110001010010111011010" OR uut_h_1_1 /= "000000001110100001011100000" OR uut_h_1_2 /= "000000010010001001111000001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0101011";
              state <= "1100111";
            ELSE
              state <= "0101111";
            END IF;
            uut_rst <= '0';
          WHEN "0101111" =>
            uut_h_0_0_i <= "000000000100111010010000010";
            uut_h_0_1_i <= "111111110010011100100011000";
            uut_h_0_2_i <= "000000000010101110010010001";
            uut_h_1_0_i <= "000000001110111011100011000";
            uut_h_1_1_i <= "000000001001010100110100010";
            uut_h_1_2_i <= "111111110101110111011110010";
            uut_xb <= "111111110100111010101100111";
            uut_yb <= "000000001010011101011100010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000011011001110100010" OR uut_h_0_1 /= "111111111111101001100011010" OR uut_h_0_2 /= "000000010011110010100010001" OR uut_h_1_0 /= "000000001010001000100101111" OR uut_h_1_1 /= "000000001000010101111110001" OR uut_h_1_2 /= "111111101100011001111110011" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0101100";
              state <= "1100111";
            ELSE
              state <= "0110000";
            END IF;
            uut_rst <= '0';
          WHEN "0110000" =>
            uut_h_0_0_i <= "111111111001101000010111000";
            uut_h_0_1_i <= "000000001010001001111110011";
            uut_h_0_2_i <= "111111110110000100110101101";
            uut_h_1_0_i <= "111111111100010010001100100";
            uut_h_1_1_i <= "000000001000100001010100000";
            uut_h_1_2_i <= "000000000100101100000010010";
            uut_xb <= "111111111001000011010110101";
            uut_yb <= "000000000100011011110110101";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000111111001101000010" OR uut_h_0_1 /= "111111111000010101100110100" OR uut_h_0_2 /= "000000010101110001110111000" OR uut_h_1_0 /= "111111111111001101111100010" OR uut_h_1_1 /= "111111110010101101101101110" OR uut_h_1_2 /= "000000001111011010001101001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0101101";
              state <= "1100111";
            ELSE
              state <= "0110001";
            END IF;
            uut_rst <= '0';
          WHEN "0110001" =>
            uut_h_0_0_i <= "000000000010111100100100011";
            uut_h_0_1_i <= "111111110011111100011000110";
            uut_h_0_2_i <= "111111111101111010001010000";
            uut_h_1_0_i <= "111111111010011010001100010";
            uut_h_1_1_i <= "000000000111100011000100110";
            uut_h_1_2_i <= "000000001010101000011011110";
            uut_xb <= "111111110010011100001000101";
            uut_yb <= "000000000001110100100101010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110000101011100111110" OR uut_h_0_1 /= "111111111010010111111000111" OR uut_h_0_2 /= "000000011100110110111000100" OR uut_h_1_0 /= "000000001100001010001101100" OR uut_h_1_1 /= "000000000101011010001100111" OR uut_h_1_2 /= "111111110010100100111000001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0101110";
              state <= "1100111";
            ELSE
              state <= "0110010";
            END IF;
            uut_rst <= '0';
          WHEN "0110010" =>
            uut_h_0_0_i <= "111111111000110001000000100";
            uut_h_0_1_i <= "111111111111100011001000100";
            uut_h_0_2_i <= "111111110110011100110110000";
            uut_h_1_0_i <= "111111110100001110011100101";
            uut_h_1_1_i <= "111111110101110110001100111";
            uut_h_1_2_i <= "111111110100010011111101011";
            uut_xb <= "000000001110011010101101110";
            uut_yb <= "000000000001000001110011011";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000100111010010000010" OR uut_h_0_1 /= "111111110010011100100011000" OR uut_h_0_2 /= "000000000011111001110000101" OR uut_h_1_0 /= "000000001110111011100011000" OR uut_h_1_1 /= "000000001001010100110100010" OR uut_h_1_2 /= "000000000100100100101000011" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0101111";
              state <= "1100111";
            ELSE
              state <= "0110011";
            END IF;
            uut_rst <= '0';
          WHEN "0110011" =>
            uut_h_0_0_i <= "111111110111111011010000101";
            uut_h_0_1_i <= "000000000001100001101011100";
            uut_h_0_2_i <= "111111111100001011101010100";
            uut_h_1_0_i <= "111111111101111111100010101";
            uut_h_1_1_i <= "000000000011011111010101111";
            uut_h_1_2_i <= "000000000111111101110111000";
            uut_xb <= "111111110001110111000010011";
            uut_yb <= "111111111010110111101110000";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111001101000010111000" OR uut_h_0_1 /= "000000001010001001111110011" OR uut_h_0_2 /= "111111101001100011000000111" OR uut_h_1_0 /= "111111111100010010001100100" OR uut_h_1_1 /= "000000001000100001010100000" OR uut_h_1_2 /= "000000000101001001011110000" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0110000";
              state <= "1100111";
            ELSE
              state <= "0110100";
            END IF;
            uut_rst <= '0';
          WHEN "0110100" =>
            uut_h_0_0_i <= "000000001010001001100100111";
            uut_h_0_1_i <= "000000000011010111101100010";
            uut_h_0_2_i <= "000000001100101111111110010";
            uut_h_1_0_i <= "111111111100000101001101111";
            uut_h_1_1_i <= "111111111010110100101101010";
            uut_h_1_2_i <= "000000001011001110001111110";
            uut_xb <= "111111111001001000101100011";
            uut_yb <= "000000001000111101010101001";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000010111100100100011" OR uut_h_0_1 /= "111111110011111100011000110" OR uut_h_0_2 /= "111111110100001101111101010" OR uut_h_1_0 /= "111111111010011010001100010" OR uut_h_1_1 /= "000000000111100011000100110" OR uut_h_1_2 /= "000000000110110110110001010" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0110001";
              state <= "1100111";
            ELSE
              state <= "0110101";
            END IF;
            uut_rst <= '0';
          WHEN "0110101" =>
            uut_h_0_0_i <= "000000000110011100011101010";
            uut_h_0_1_i <= "111111111111001111001011011";
            uut_h_0_2_i <= "000000000000000111000100101";
            uut_h_1_0_i <= "111111111111110000101010100";
            uut_h_1_1_i <= "000000001111110101100100010";
            uut_h_1_2_i <= "000000001000100110011100100";
            uut_xb <= "111111111110100000010001100";
            uut_yb <= "111111110100010000000101011";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111000110001000000100" OR uut_h_0_1 /= "111111111111100011001000100" OR uut_h_0_2 /= "000000001011011010100111001" OR uut_h_1_0 /= "111111110100001110011100101" OR uut_h_1_1 /= "111111110101110110001100111" OR uut_h_1_2 /= "000000000000100110100010100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0110010";
              state <= "1100111";
            ELSE
              state <= "0110110";
            END IF;
            uut_rst <= '0';
          WHEN "0110110" =>
            uut_h_0_0_i <= "000000001000010001011010111";
            uut_h_0_1_i <= "000000001001100010011011000";
            uut_h_0_2_i <= "000000001100111100111000101";
            uut_h_1_0_i <= "000000000010000101100110101";
            uut_h_1_1_i <= "111111110111000011011110100";
            uut_h_1_2_i <= "111111111001010110000011101";
            uut_xb <= "111111111010110111001011110";
            uut_yb <= "111111111000101110011100110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110111111011010000101" OR uut_h_0_1 /= "000000000001100001101011100" OR uut_h_0_2 /= "111111100111011001010110010" OR uut_h_1_0 /= "111111111101111111100010101" OR uut_h_1_1 /= "000000000011011111010101111" OR uut_h_1_2 /= "000000000010001011101001111" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0110011";
              state <= "1100111";
            ELSE
              state <= "0110111";
            END IF;
            uut_rst <= '0';
          WHEN "0110111" =>
            uut_h_0_0_i <= "111111110101011100101110001";
            uut_h_0_1_i <= "000000001010100010000001000";
            uut_h_0_2_i <= "111111111101110011000100011";
            uut_h_1_0_i <= "000000000101001111111010001";
            uut_h_1_1_i <= "111111111000100011100011101";
            uut_h_1_2_i <= "111111111111001110001001000";
            uut_xb <= "111111110100001011100100110";
            uut_yb <= "111111110001101001001011010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001010001001100100111" OR uut_h_0_1 /= "000000000011010111101100010" OR uut_h_0_2 /= "000000001000010110100101000" OR uut_h_1_0 /= "111111111100000101001101111" OR uut_h_1_1 /= "111111111010110100101101010" OR uut_h_1_2 /= "000000010101011001011110101" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0110100";
              state <= "1100111";
            ELSE
              state <= "0111000";
            END IF;
            uut_rst <= '0';
          WHEN "0111000" =>
            uut_h_0_0_i <= "000000000100000101001000100";
            uut_h_0_1_i <= "000000000110001110011100110";
            uut_h_0_2_i <= "000000001001110111110001100";
            uut_h_1_0_i <= "111111110000111011100100100";
            uut_h_1_1_i <= "000000000000100000000111000";
            uut_h_1_2_i <= "000000001001011001011110000";
            uut_xb <= "111111111000110110100010101";
            uut_yb <= "111111110011110101000100101";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000110011100011101010" OR uut_h_0_1 /= "111111111111001111001011011" OR uut_h_0_2 /= "111111111110101010000011100" OR uut_h_1_0 /= "111111111111110000101010100" OR uut_h_1_1 /= "000000001111110101100100010" OR uut_h_1_2 /= "000000001000011101010110100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0110101";
              state <= "1100111";
            ELSE
              state <= "0111001";
            END IF;
            uut_rst <= '0';
          WHEN "0111001" =>
            uut_h_0_0_i <= "000000001100010111110000001";
            uut_h_0_1_i <= "000000000100011010111000101";
            uut_h_0_2_i <= "111111110101110101101010001";
            uut_h_1_0_i <= "000000001111000011001001101";
            uut_h_1_1_i <= "111111110010111001100001110";
            uut_h_1_2_i <= "111111110001000000111001010";
            uut_xb <= "111111110100100111001111001";
            uut_yb <= "000000000100010110011000001";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001000010001011010111" OR uut_h_0_1 /= "000000001001100010011011000" OR uut_h_0_2 /= "000000001110110011100110000" OR uut_h_1_0 /= "000000000010000101100110101" OR uut_h_1_1 /= "111111110111000011011110100" OR uut_h_1_2 /= "111111101110101011000111100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0110110";
              state <= "1100111";
            ELSE
              state <= "0111010";
            END IF;
            uut_rst <= '0';
          WHEN "0111010" =>
            uut_h_0_0_i <= "000000001001010001100110111";
            uut_h_0_1_i <= "000000001010010010100110111";
            uut_h_0_2_i <= "000000001001000111101000111";
            uut_h_1_0_i <= "000000000010000111101011111";
            uut_h_1_1_i <= "111111111001110000011001010";
            uut_h_1_2_i <= "000000000000000111101001101";
            uut_xb <= "000000000111011100000111000";
            uut_yb <= "111111110101001101101110001";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110101011100101110001" OR uut_h_0_1 /= "000000001010100010000001000" OR uut_h_0_2 /= "111111110011101000100110101" OR uut_h_1_0 /= "000000000101001111111010001" OR uut_h_1_1 /= "111111111000100011100011101" OR uut_h_1_2 /= "111111101110000011111100100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0110111";
              state <= "1100111";
            ELSE
              state <= "0111011";
            END IF;
            uut_rst <= '0';
          WHEN "0111011" =>
            uut_h_0_0_i <= "000000001101011110010111001";
            uut_h_0_1_i <= "111111110010010110111100001";
            uut_h_0_2_i <= "000000000111101100011001000";
            uut_h_1_0_i <= "111111110111000111000111010";
            uut_h_1_1_i <= "000000001000101000000010101";
            uut_h_1_2_i <= "000000001000010000111001001";
            uut_xb <= "111111111110111011001111010";
            uut_yb <= "000000001001001011110001001";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000100000101001000100" OR uut_h_0_1 /= "000000000110001110011100110" OR uut_h_0_2 /= "000000001001010010000100000" OR uut_h_1_0 /= "111111110000111011100100100" OR uut_h_1_1 /= "000000000000100000000111000" OR uut_h_1_2 /= "111111110110111000000111110" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0111000";
              state <= "1100111";
            ELSE
              state <= "0111100";
            END IF;
            uut_rst <= '0';
          WHEN "0111100" =>
            uut_h_0_0_i <= "111111111101100001011010110";
            uut_h_0_1_i <= "000000001111011001101000101";
            uut_h_0_2_i <= "000000000001110101110001000";
            uut_h_1_0_i <= "000000001110001100110000100";
            uut_h_1_1_i <= "000000000010001111110000011";
            uut_h_1_2_i <= "111111111001100101111101011";
            uut_xb <= "000000000101010010011100011";
            uut_yb <= "000000000101111001001111110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001100010111110000001" OR uut_h_0_1 /= "000000000100011010111000101" OR uut_h_0_2 /= "111111110010000011011110001" OR uut_h_1_0 /= "000000001111000011001001101" OR uut_h_1_1 /= "111111110010111001100001110" OR uut_h_1_2 /= "000000000011101000101011000" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0111001";
              state <= "1100111";
            ELSE
              state <= "0111101";
            END IF;
            uut_rst <= '0';
          WHEN "0111101" =>
            uut_h_0_0_i <= "000000001001010110110110101";
            uut_h_0_1_i <= "111111111011000010100100010";
            uut_h_0_2_i <= "000000001000001100011011111";
            uut_h_1_0_i <= "111111111011001001111110111";
            uut_h_1_1_i <= "111111111010100001000010100";
            uut_h_1_2_i <= "111111111001001110010100000";
            uut_xb <= "000000001000100000110101000";
            uut_yb <= "000000001011000100111010111";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001001010001100110111" OR uut_h_0_1 /= "000000001010010010100110111" OR uut_h_0_2 /= "000000010011001011101110000" OR uut_h_1_0 /= "000000000010000111101011111" OR uut_h_1_1 /= "111111111001110000011001010" OR uut_h_1_2 /= "111111110000001000111010011" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0111010";
              state <= "1100111";
            ELSE
              state <= "0111110";
            END IF;
            uut_rst <= '0';
          WHEN "0111110" =>
            uut_h_0_0_i <= "000000001100110111010000011";
            uut_h_0_1_i <= "111111110110111110100011011";
            uut_h_0_2_i <= "000000000101001010001010000";
            uut_h_1_0_i <= "000000000011000100000000100";
            uut_h_1_1_i <= "000000001011110100100011000";
            uut_h_1_2_i <= "000000001001000100100100111";
            uut_xb <= "000000000001101111011101101";
            uut_yb <= "111111110111010110001100001";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001101011110010111001" OR uut_h_0_1 /= "111111110010010110111100001" OR uut_h_0_2 /= "000000001111010110101010110" OR uut_h_1_0 /= "111111110111000111000111010" OR uut_h_1_1 /= "000000001000101000000010101" OR uut_h_1_2 /= "000000001011111001100110001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0111011";
              state <= "1100111";
            ELSE
              state <= "0111111";
            END IF;
            uut_rst <= '0';
          WHEN "0111111" =>
            uut_h_0_0_i <= "111111110000001110001010000";
            uut_h_0_1_i <= "111111111100100101000100110";
            uut_h_0_2_i <= "000000000101001100010110010";
            uut_h_1_0_i <= "000000001000100010000100111";
            uut_h_1_1_i <= "111111111000000101001100111";
            uut_h_1_2_i <= "000000001101010001011001000";
            uut_xb <= "000000000111111000101011001";
            uut_yb <= "000000001001100101101110011";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111101100001011010110" OR uut_h_0_1 /= "000000001111011001101000101" OR uut_h_0_2 /= "000000000010010001100000110" OR uut_h_1_0 /= "000000001110001100110000100" OR uut_h_1_1 /= "000000000010001111110000011" OR uut_h_1_2 /= "111111111001111101111001001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0111100";
              state <= "1100111";
            ELSE
              state <= "1000000";
            END IF;
            uut_rst <= '0';
          WHEN "1000000" =>
            uut_h_0_0_i <= "000000001101000011001011000";
            uut_h_0_1_i <= "000000000000100110110110011";
            uut_h_0_2_i <= "000000001110100001100110111";
            uut_h_1_0_i <= "000000001111001011111011010";
            uut_h_1_1_i <= "000000001010010011011001111";
            uut_h_1_2_i <= "000000001110010011010011100";
            uut_xb <= "111111110010001001111010111";
            uut_yb <= "111111111110000000000100100";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001001010110110110101" OR uut_h_0_1 /= "111111111011000010100100010" OR uut_h_0_2 /= "000000001111001010011001101" OR uut_h_1_0 /= "111111111011001001111110111" OR uut_h_1_1 /= "111111111010100001000010100" OR uut_h_1_2 /= "000000001010101011001001111" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0111101";
              state <= "1100111";
            ELSE
              state <= "1000001";
            END IF;
            uut_rst <= '0';
          WHEN "1000001" =>
            uut_h_0_0_i <= "111111111010010001000101001";
            uut_h_0_1_i <= "000000001001110010100101001";
            uut_h_0_2_i <= "000000001111101000000111101";
            uut_h_1_0_i <= "111111110100010010100010011";
            uut_h_1_1_i <= "000000000000110010101101111";
            uut_h_1_2_i <= "111111111101000111011101101";
            uut_xb <= "111111110111010000100110001";
            uut_yb <= "111111111110010001011110001";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001100110111010000011" OR uut_h_0_1 /= "111111110110111110100011011" OR uut_h_0_2 /= "000000000000100111101101010" OR uut_h_1_0 /= "000000000011000100000000100" OR uut_h_1_1 /= "000000001011110100100011000" OR uut_h_1_2 /= "000000000110011110100110001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0111110";
              state <= "1100111";
            ELSE
              state <= "1000010";
            END IF;
            uut_rst <= '0';
          WHEN "1000010" =>
            uut_h_0_0_i <= "111111111000100001001110001";
            uut_h_0_1_i <= "111111111000010011101101010";
            uut_h_0_2_i <= "000000000000001110000011001";
            uut_h_1_0_i <= "111111111110101100001110101";
            uut_h_1_1_i <= "111111110100010001110110001";
            uut_h_1_2_i <= "111111111010011000001101110";
            uut_xb <= "111111111110001011011101001";
            uut_yb <= "111111111101111100001111001";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110000001110001010000" OR uut_h_0_1 /= "111111111100100101000100110" OR uut_h_0_2 /= "000000010110111001111011101" OR uut_h_1_0 /= "000000001000100010000100111" OR uut_h_1_1 /= "111111111000000101001100111" OR uut_h_1_2 /= "000000010111011001101110110" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "0111111";
              state <= "1100111";
            ELSE
              state <= "1000011";
            END IF;
            uut_rst <= '0';
          WHEN "1000011" =>
            uut_h_0_0_i <= "000000001001011000000111001";
            uut_h_0_1_i <= "000000001001010000011001010";
            uut_h_0_2_i <= "000000000100001011110001101";
            uut_h_1_0_i <= "000000001010000110010000100";
            uut_h_1_1_i <= "000000000000000010100110001";
            uut_h_1_2_i <= "111111110011001000101011101";
            uut_xb <= "000000000011101101000000010";
            uut_yb <= "111111111001110000100011101";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001101000011001011000" OR uut_h_0_1 /= "000000000000100110110110011" OR uut_h_0_2 /= "000000001100000011000100011" OR uut_h_1_0 /= "000000001111001011111011010" OR uut_h_1_1 /= "000000001010010011011001111" OR uut_h_1_2 /= "000000011010101110110001110" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1000000";
              state <= "1100111";
            ELSE
              state <= "1000100";
            END IF;
            uut_rst <= '0';
          WHEN "1000100" =>
            uut_h_0_0_i <= "000000001000100010101111111";
            uut_h_0_1_i <= "111111111001011111010110111";
            uut_h_0_2_i <= "000000000110000011010100111";
            uut_h_1_0_i <= "111111111000100011010010010";
            uut_h_1_1_i <= "000000000001110011011011110";
            uut_h_1_2_i <= "000000000110111110001110001";
            uut_xb <= "000000000001000100010011110";
            uut_yb <= "000000001100000001011110111";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111010010001000101001" OR uut_h_0_1 /= "000000001001110010100101001" OR uut_h_0_2 /= "000000000100110011111001110" OR uut_h_1_0 /= "111111110100010010100010011" OR uut_h_1_1 /= "000000000000110010101101111" OR uut_h_1_2 /= "111111110101000100111110111" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1000001";
              state <= "1100111";
            ELSE
              state <= "1000101";
            END IF;
            uut_rst <= '0';
          WHEN "1000101" =>
            uut_h_0_0_i <= "111111111100100101000100001";
            uut_h_0_1_i <= "000000001000001110111001010";
            uut_h_0_2_i <= "000000000110011011101001001";
            uut_h_1_0_i <= "111111111110101010000111101";
            uut_h_1_1_i <= "000000000001011111101000000";
            uut_h_1_2_i <= "111111110011011111101100000";
            uut_xb <= "000000000011000111010001100";
            uut_yb <= "000000000101000101111111100";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111000100001001110001" OR uut_h_0_1 /= "111111111000010011101101010" OR uut_h_0_2 /= "111111111100100011101010110" OR uut_h_1_0 /= "111111111110101100001110101" OR uut_h_1_1 /= "111111110100010001110110001" OR uut_h_1_2 /= "111111110110101010011001001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1000010";
              state <= "1100111";
            ELSE
              state <= "1000110";
            END IF;
            uut_rst <= '0';
          WHEN "1000110" =>
            uut_h_0_0_i <= "000000000010100011110110100";
            uut_h_0_1_i <= "000000000000110100010110010";
            uut_h_0_2_i <= "000000000111011011000010001";
            uut_h_1_0_i <= "000000001101000111100101001";
            uut_h_1_1_i <= "111111111000010011101101010";
            uut_h_1_2_i <= "111111110101010000011110000";
            uut_xb <= "111111111000010011010011101";
            uut_yb <= "000000000001100000011100111";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001001011000000111001" OR uut_h_0_1 /= "000000001001010000011001010" OR uut_h_0_2 /= "000000001001010100111110000" OR uut_h_1_0 /= "000000001010000110010000100" OR uut_h_1_1 /= "000000000000000010100110001" OR uut_h_1_2 /= "111111101010100100101011011" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1000011";
              state <= "1100111";
            ELSE
              state <= "1000111";
            END IF;
            uut_rst <= '0';
          WHEN "1000111" =>
            uut_h_0_0_i <= "000000000001010100100001001";
            uut_h_0_1_i <= "000000001001001100111000100";
            uut_h_0_2_i <= "000000001101110001110111011";
            uut_h_1_0_i <= "000000001001001110000011100";
            uut_h_1_1_i <= "000000001111000001011000110";
            uut_h_1_2_i <= "111111110001011100011110001";
            uut_xb <= "111111110000010010001000101";
            uut_yb <= "000000000101011111011011000";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001000100010101111111" OR uut_h_0_1 /= "111111111001011111010110111" OR uut_h_0_2 /= "000000001011011100010000000" OR uut_h_1_0 /= "111111111000100011010010010" OR uut_h_1_1 /= "000000000001110011011011110" OR uut_h_1_2 /= "000000010010001000110000110" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1000100";
              state <= "1100111";
            ELSE
              state <= "1001000";
            END IF;
            uut_rst <= '0';
          WHEN "1001000" =>
            uut_h_0_0_i <= "000000001100111101000011101";
            uut_h_0_1_i <= "000000000000000100110110010";
            uut_h_0_2_i <= "111111111010010111111101000";
            uut_h_1_0_i <= "000000000010010100010011110";
            uut_h_1_1_i <= "000000000010001010101101111";
            uut_h_1_2_i <= "000000000110111010011100011";
            uut_xb <= "111111110100100011011001001";
            uut_yb <= "111111111100001010111111000";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111100100101000100001" OR uut_h_0_1 /= "000000001000001110111001010" OR uut_h_0_2 /= "000000000111100101110010011" OR uut_h_1_0 /= "111111111110101010000111101" OR uut_h_1_1 /= "000000000001011111101000000" OR uut_h_1_2 /= "111111111000010111111100111" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1000101";
              state <= "1100111";
            ELSE
              state <= "1001001";
            END IF;
            uut_rst <= '0';
          WHEN "1001001" =>
            uut_h_0_0_i <= "111111111100101100001011000";
            uut_h_0_1_i <= "000000000010011110111000100";
            uut_h_0_2_i <= "000000000111011011011100010";
            uut_h_1_0_i <= "000000000010011101001010101";
            uut_h_1_1_i <= "000000001101110101001000110";
            uut_h_1_2_i <= "000000001111000011101000010";
            uut_xb <= "000000000111000001111000000";
            uut_yb <= "111111111001101100000010010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000010100011110110100" OR uut_h_0_1 /= "000000000000110100010110010" OR uut_h_0_2 /= "000000000000111000001111111" OR uut_h_1_0 /= "000000001101000111100101001" OR uut_h_1_1 /= "111111111000010011101101010" OR uut_h_1_2 /= "111111111101110011010000001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1000110";
              state <= "1100111";
            ELSE
              state <= "1001010";
            END IF;
            uut_rst <= '0';
          WHEN "1001010" =>
            uut_h_0_0_i <= "111111111110101100000100111";
            uut_h_0_1_i <= "111111111011100100110010111";
            uut_h_0_2_i <= "111111111110011010101011100";
            uut_h_1_0_i <= "111111110001100010010111001";
            uut_h_1_1_i <= "111111111001001100111110001";
            uut_h_1_2_i <= "000000001001110011111110111";
            uut_xb <= "111111111001000011011111110";
            uut_yb <= "111111110010001011111001011";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000001010100100001001" OR uut_h_0_1 /= "000000001001001100111000100" OR uut_h_0_2 /= "111111111100001100111011010" OR uut_h_1_0 /= "000000001001001110000011100" OR uut_h_1_1 /= "000000001111000001011000110" OR uut_h_1_2 /= "111111111010110101100100001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1000111";
              state <= "1100111";
            ELSE
              state <= "1001011";
            END IF;
            uut_rst <= '0';
          WHEN "1001011" =>
            uut_h_0_0_i <= "111111110001110000011111111";
            uut_h_0_1_i <= "000000001100111110100001110";
            uut_h_0_2_i <= "000000000001010001111010110";
            uut_h_1_0_i <= "000000000100011001101001010";
            uut_h_1_1_i <= "111111111101010110101011000";
            uut_h_1_2_i <= "000000001101111111001010011";
            uut_xb <= "111111111100101000010000100";
            uut_yb <= "111111111000010010011010011";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001100111101000011101" OR uut_h_0_1 /= "000000000000000100110110010" OR uut_h_0_2 /= "111111111000001101101001010" OR uut_h_1_0 /= "000000000010010100010011110" OR uut_h_1_1 /= "000000000010001010101101111" OR uut_h_1_2 /= "000000000101010000101110011" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1001000";
              state <= "1100111";
            ELSE
              state <= "1001100";
            END IF;
            uut_rst <= '0';
          WHEN "1001100" =>
            uut_h_0_0_i <= "000000001011001000100001100";
            uut_h_0_1_i <= "111111110010001001110010100";
            uut_h_0_2_i <= "111111110101111100101100010";
            uut_h_1_0_i <= "000000001110001111011110011";
            uut_h_1_1_i <= "111111110101110011111000010";
            uut_h_1_2_i <= "111111111001010100111000101";
            uut_xb <= "111111111011000110100111000";
            uut_yb <= "111111111010001011100110100";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111100101100001011000" OR uut_h_0_1 /= "000000000010011110111000100" OR uut_h_0_2 /= "000000010000111001000011111" OR uut_h_1_0 /= "000000000010011101001010101" OR uut_h_1_1 /= "000000001101110101001000110" OR uut_h_1_2 /= "000000001101000111110011011" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1001001";
              state <= "1100111";
            ELSE
              state <= "1001101";
            END IF;
            uut_rst <= '0';
          WHEN "1001101" =>
            uut_h_0_0_i <= "111111111110101101111001111";
            uut_h_0_1_i <= "000000000101000100100000110";
            uut_h_0_2_i <= "111111111101000100110001010";
            uut_h_1_0_i <= "111111110111100011000111001";
            uut_h_1_1_i <= "111111110101000101001110101";
            uut_h_1_2_i <= "111111111010011110011111111";
            uut_xb <= "000000000111111000100001110";
            uut_yb <= "111111110101100100010000101";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111110101100000100111" OR uut_h_0_1 /= "111111111011100100110010111" OR uut_h_0_2 /= "111111110011000101001110111" OR uut_h_1_0 /= "111111110001100010010111001" OR uut_h_1_1 /= "111111111001001100111110001" OR uut_h_1_2 /= "111111101111110110011110100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1001010";
              state <= "1100111";
            ELSE
              state <= "1001110";
            END IF;
            uut_rst <= '0';
          WHEN "1001110" =>
            uut_h_0_0_i <= "111111110011110000101110110";
            uut_h_0_1_i <= "000000001010111100001100001";
            uut_h_0_2_i <= "000000000110110110111001011";
            uut_h_1_0_i <= "111111110101100100011011011";
            uut_h_1_1_i <= "000000000000010100101001100";
            uut_h_1_2_i <= "000000001101000001100111001";
            uut_xb <= "000000001011110111101110101";
            uut_yb <= "111111110110110001110101110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110001110000011111111" OR uut_h_0_1 /= "000000001100111110100001110" OR uut_h_0_2 /= "000000000001001010011110000" OR uut_h_1_0 /= "000000000100011001101001010" OR uut_h_1_1 /= "111111111101010110101011000" OR uut_h_1_2 /= "000000000101111011010010111" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1001011";
              state <= "1100111";
            ELSE
              state <= "1001111";
            END IF;
            uut_rst <= '0';
          WHEN "1001111" =>
            uut_h_0_0_i <= "000000001010110001011111010";
            uut_h_0_1_i <= "111111111111010001101000111";
            uut_h_0_2_i <= "000000000000010011010111011";
            uut_h_1_0_i <= "000000001011011111110110011";
            uut_h_1_1_i <= "000000001100011110011110110";
            uut_h_1_2_i <= "000000000011110111011001001";
            uut_xb <= "111111110111010111000010000";
            uut_yb <= "111111110000101100110010110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001011001000100001100" OR uut_h_0_1 /= "111111110010001001110010100" OR uut_h_0_2 /= "111111101111011011000101001" OR uut_h_1_0 /= "000000001110001111011110011" OR uut_h_1_1 /= "111111110101110011111000010" OR uut_h_1_2 /= "111111110100001010010010001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1001100";
              state <= "1100111";
            ELSE
              state <= "1010000";
            END IF;
            uut_rst <= '0';
          WHEN "1010000" =>
            uut_h_0_0_i <= "111111110100011100101001100";
            uut_h_0_1_i <= "111111111100011000001001111";
            uut_h_0_2_i <= "111111110100011000111001111";
            uut_h_1_0_i <= "000000001000100111111100111";
            uut_h_1_1_i <= "000000001111110010100010100";
            uut_h_1_2_i <= "111111111100010011111110011";
            uut_xb <= "000000000100010010000110000";
            uut_yb <= "000000000001010101001101011";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111110101101111001111" OR uut_h_0_1 /= "000000000101000100100000110" OR uut_h_0_2 /= "000000001000111001010110111" OR uut_h_1_0 /= "111111110111100011000111001" OR uut_h_1_1 /= "111111110101000101001110101" OR uut_h_1_2 /= "111111101101000101100110001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1001101";
              state <= "1100111";
            ELSE
              state <= "1010001";
            END IF;
            uut_rst <= '0';
          WHEN "1010001" =>
            uut_h_0_0_i <= "111111111010000101000110110";
            uut_h_0_1_i <= "111111110100011000011110011";
            uut_h_0_2_i <= "111111110011100111111110101";
            uut_h_1_0_i <= "111111110101000110010011010";
            uut_h_1_1_i <= "000000000110101101101011010";
            uut_h_1_2_i <= "000000000110011011011001100";
            uut_xb <= "000000001001101101111010011";
            uut_yb <= "000000000000011100100101010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110011110000101110110" OR uut_h_0_1 /= "000000001010111100001100001" OR uut_h_0_2 /= "000000100010000111010010101" OR uut_h_1_0 /= "111111110101100100011011011" OR uut_h_1_1 /= "000000000000010100101001100" OR uut_h_1_2 /= "000000001011101110101000111" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1001110";
              state <= "1100111";
            ELSE
              state <= "1010010";
            END IF;
            uut_rst <= '0';
          WHEN "1010010" =>
            uut_h_0_0_i <= "000000000001100011001100111";
            uut_h_0_1_i <= "000000000000110110010000000";
            uut_h_0_2_i <= "000000000111000100111011011";
            uut_h_1_0_i <= "111111110110101001101010101";
            uut_h_1_1_i <= "000000000010010001011101001";
            uut_h_1_2_i <= "111111110010010101110010011";
            uut_xb <= "000000001011100101010101000";
            uut_yb <= "111111111110010111001001010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001010110001011111010" OR uut_h_0_1 /= "111111111111010001101000111" OR uut_h_0_2 /= "111111111100110010011001010" OR uut_h_1_0 /= "000000001011011111110110011" OR uut_h_1_1 /= "000000001100011110011110110" OR uut_h_1_2 /= "000000000110101101000110101" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1001111";
              state <= "1100111";
            ELSE
              state <= "1010011";
            END IF;
            uut_rst <= '0';
          WHEN "1010011" =>
            uut_h_0_0_i <= "000000000100111000011110100";
            uut_h_0_1_i <= "111111111000111011001100010";
            uut_h_0_2_i <= "000000001110100001111110000";
            uut_h_1_0_i <= "111111111001101101100000110";
            uut_h_1_1_i <= "000000001001100101100000001";
            uut_h_1_2_i <= "111111111110001110000000010";
            uut_xb <= "000000000011001100011011001";
            uut_yb <= "000000001010111101101100001";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110100011100101001100" OR uut_h_0_1 /= "111111111100011000001001111" OR uut_h_0_2 /= "111111111100000100001100011" OR uut_h_1_0 /= "000000001000100111111100111" OR uut_h_1_1 /= "000000001111110010100010100" OR uut_h_1_2 /= "111111111010000001010110110" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1010000";
              state <= "1100111";
            ELSE
              state <= "1010100";
            END IF;
            uut_rst <= '0';
          WHEN "1010100" =>
            uut_h_0_0_i <= "111111110000111111111001100";
            uut_h_0_1_i <= "000000001110010101010110000";
            uut_h_0_2_i <= "000000001101101110010110000";
            uut_h_1_0_i <= "111111110101111111100001110";
            uut_h_1_1_i <= "111111111110011111101101100";
            uut_h_1_2_i <= "000000000101100001101110011";
            uut_xb <= "111111111100111110110111010";
            uut_yb <= "111111111110000010101101100";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111010000101000110110" OR uut_h_0_1 /= "111111110100011000011110011" OR uut_h_0_2 /= "000000000001010000110000110" OR uut_h_1_0 /= "111111110101000110010011010" OR uut_h_1_1 /= "000000000110101101101011010" OR uut_h_1_2 /= "000000001101010011101110100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1010001";
              state <= "1100111";
            ELSE
              state <= "1010101";
            END IF;
            uut_rst <= '0';
          WHEN "1010101" =>
            uut_h_0_0_i <= "000000000101101101110111111";
            uut_h_0_1_i <= "111111111011010110011010111";
            uut_h_0_2_i <= "000000000001011101000011001";
            uut_h_1_0_i <= "111111111110111000011101101";
            uut_h_1_1_i <= "111111111010110110010100001";
            uut_h_1_2_i <= "000000000111111110100010000";
            uut_xb <= "111111111110100000001110011";
            uut_yb <= "111111110010011001000101100";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000001100011001100111" OR uut_h_0_1 /= "000000000000110110010000000" OR uut_h_0_2 /= "000000010001100111111111110" OR uut_h_1_0 /= "111111110110101001101010101" OR uut_h_1_1 /= "000000000010010001011101001" OR uut_h_1_2 /= "111111110111101100111111100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1010010";
              state <= "1100111";
            ELSE
              state <= "1010110";
            END IF;
            uut_rst <= '0';
          WHEN "1010110" =>
            uut_h_0_0_i <= "000000000101001110100001011";
            uut_h_0_1_i <= "000000000101000111110100111";
            uut_h_0_2_i <= "111111111110111110010000110";
            uut_h_1_0_i <= "000000000110100001000101000";
            uut_h_1_1_i <= "000000000110000101010101011";
            uut_h_1_2_i <= "111111111110101010111101101";
            uut_xb <= "000000001010011001000111111";
            uut_yb <= "111111110110000110000000110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000100111000011110100" OR uut_h_0_1 /= "111111111000111011001100010" OR uut_h_0_2 /= "000000010101100110010011001" OR uut_h_1_0 /= "111111111001101101100000110" OR uut_h_1_1 /= "000000001001100101100000001" OR uut_h_1_2 /= "000000000011110111101001100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1010011";
              state <= "1100111";
            ELSE
              state <= "1010111";
            END IF;
            uut_rst <= '0';
          WHEN "1010111" =>
            uut_h_0_0_i <= "111111110000110100100101000";
            uut_h_0_1_i <= "111111110101011111000100001";
            uut_h_0_2_i <= "111111111111000111010101100";
            uut_h_1_0_i <= "111111110001110100010110110";
            uut_h_1_1_i <= "000000000100000001101110101";
            uut_h_1_2_i <= "000000000101101101011100110";
            uut_xb <= "111111110111100011011101010";
            uut_yb <= "111111111001010000000010010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110000111111111001100" OR uut_h_0_1 /= "000000001110010101010110000" OR uut_h_0_2 /= "000000001001101000010111010" OR uut_h_1_0 /= "111111110101111111100001110" OR uut_h_1_1 /= "111111111110011111101101100" OR uut_h_1_2 /= "000000000001011111110110111" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1010100";
              state <= "1100111";
            ELSE
              state <= "1011000";
            END IF;
            uut_rst <= '0';
          WHEN "1011000" =>
            uut_h_0_0_i <= "111111110101100001110011100";
            uut_h_0_1_i <= "111111111001100101101001100";
            uut_h_0_2_i <= "000000000001110000000000100";
            uut_h_1_0_i <= "111111111010010110111100110";
            uut_h_1_1_i <= "000000001000110100011110110";
            uut_h_1_2_i <= "000000000111011000010111011";
            uut_xb <= "000000001100110100111011110";
            uut_yb <= "111111110100011010111101110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000101101101110111111" OR uut_h_0_1 /= "111111111011010110011010111" OR uut_h_0_2 /= "111111111100100010011001110" OR uut_h_1_0 /= "111111111110111000011101101" OR uut_h_1_1 /= "111111111010110110010100001" OR uut_h_1_2 /= "111111110101111000100010000" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1010101";
              state <= "1100111";
            ELSE
              state <= "1011001";
            END IF;
            uut_rst <= '0';
          WHEN "1011001" =>
            uut_h_0_0_i <= "000000001001011010010001001";
            uut_h_0_1_i <= "111111110100000100111000111";
            uut_h_0_2_i <= "000000001101111011011010010";
            uut_h_1_0_i <= "111111110110000011111010110";
            uut_h_1_1_i <= "111111110100010001111001000";
            uut_h_1_2_i <= "111111111000101111100100110";
            uut_xb <= "000000000100011010111011101";
            uut_yb <= "000000001011111010111100010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000101001110100001011" OR uut_h_0_1 /= "000000000101000111110100111" OR uut_h_0_2 /= "000000001001001001000100100" OR uut_h_1_0 /= "000000000110100001000101000" OR uut_h_1_1 /= "000000000110000101010101011" OR uut_h_1_2 /= "111111110100010011000111100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1010110";
              state <= "1100111";
            ELSE
              state <= "1011010";
            END IF;
            uut_rst <= '0';
          WHEN "1011010" =>
            uut_h_0_0_i <= "111111111011101111110001000";
            uut_h_0_1_i <= "000000000001011101011111010";
            uut_h_0_2_i <= "111111110000011111110101111";
            uut_h_1_0_i <= "111111110111100011101111011";
            uut_h_1_1_i <= "111111111000001010011110100";
            uut_h_1_2_i <= "000000000010110011001011001";
            uut_xb <= "000000001011001100011111001";
            uut_yb <= "111111110000010000010000110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110000110100100101000" OR uut_h_0_1 /= "111111110101011111000100001" OR uut_h_0_2 /= "111111101010001110001000101" OR uut_h_1_0 /= "111111110001110100010110110" OR uut_h_1_1 /= "000000000100000001101110101" OR uut_h_1_2 /= "111111111001001011000101011" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1010111";
              state <= "1100111";
            ELSE
              state <= "1011011";
            END IF;
            uut_rst <= '0';
          WHEN "1011011" =>
            uut_h_0_0_i <= "000000000100010010011110111";
            uut_h_0_1_i <= "000000000001010011100110000";
            uut_h_0_2_i <= "000000001100010110110001111";
            uut_h_1_0_i <= "111111111011011111110101000";
            uut_h_1_1_i <= "111111111101010100110101001";
            uut_h_1_2_i <= "111111110100110001111101100";
            uut_xb <= "111111110001111000111010010";
            uut_yb <= "111111111100001100010110010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110101100001110011100" OR uut_h_0_1 /= "111111111001100101101001100" OR uut_h_0_2 /= "000000010010010101010001101" OR uut_h_1_0 /= "111111111010010110111100110" OR uut_h_1_1 /= "000000001000110100011110110" OR uut_h_1_2 /= "000000000110101101010001111" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1011000";
              state <= "1100111";
            ELSE
              state <= "1011100";
            END IF;
            uut_rst <= '0';
          WHEN "1011100" =>
            uut_h_0_0_i <= "000000000111000111011010011";
            uut_h_0_1_i <= "111111111001011111000001110";
            uut_h_0_2_i <= "111111111101111101101100110";
            uut_h_1_0_i <= "111111110011000010110011011";
            uut_h_1_1_i <= "000000000011001001110110110";
            uut_h_1_2_i <= "111111110000011001111110010";
            uut_xb <= "111111111000011100000001000";
            uut_yb <= "000000000000010111010100010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000001001011010010001001" OR uut_h_0_1 /= "111111110100000100111000111" OR uut_h_0_2 /= "000000011000101000100000000" OR uut_h_1_0 /= "111111110110000011111010110" OR uut_h_1_1 /= "111111110100010001111001000" OR uut_h_1_2 /= "000000010000001001001001001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1011001";
              state <= "1100111";
            ELSE
              state <= "1011101";
            END IF;
            uut_rst <= '0';
          WHEN "1011101" =>
            uut_h_0_0_i <= "111111110110111000011111100";
            uut_h_0_1_i <= "111111111101001111000101111";
            uut_h_0_2_i <= "111111111111001011101111100";
            uut_h_1_0_i <= "111111111011000100110101010";
            uut_h_1_1_i <= "111111110001110010001011100";
            uut_h_1_2_i <= "000000001010011010010000011";
            uut_xb <= "000000001010010011000001101";
            uut_yb <= "000000000010000110100000110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111011101111110001000" OR uut_h_0_1 /= "000000000001011101011111010" OR uut_h_0_2 /= "000000000000000110110100001" OR uut_h_1_0 /= "111111110111100011101111011" OR uut_h_1_1 /= "111111111000001010011110100" OR uut_h_1_2 /= "111111110001001111111001010" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1011010";
              state <= "1100111";
            ELSE
              state <= "1011110";
            END IF;
            uut_rst <= '0';
          WHEN "1011110" =>
            uut_h_0_0_i <= "111111110001101111010111111";
            uut_h_0_1_i <= "111111111111010110011111101";
            uut_h_0_2_i <= "000000001000111101110101100";
            uut_h_1_0_i <= "111111111000010100100000100";
            uut_h_1_1_i <= "111111110110010110110101100";
            uut_h_1_2_i <= "000000000011110000010000000";
            uut_xb <= "000000000110111010101000110";
            uut_yb <= "111111111100110110010010010";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000100010010011110111" OR uut_h_0_1 /= "000000000001010011100110000" OR uut_h_0_2 /= "000000000010010101101001111" OR uut_h_1_0 /= "111111111011011111110101000" OR uut_h_1_1 /= "111111111101010100110101001" OR uut_h_1_2 /= "111111101100010111011100000" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1011011";
              state <= "1100111";
            ELSE
              state <= "1011111";
            END IF;
            uut_rst <= '0';
          WHEN "1011111" =>
            uut_h_0_0_i <= "111111111110110010111101110";
            uut_h_0_1_i <= "111111110000011101011101100";
            uut_h_0_2_i <= "111111111110010001011010010";
            uut_h_1_0_i <= "000000000110101000100000110";
            uut_h_1_1_i <= "111111110010011000110111010";
            uut_h_1_2_i <= "000000001101101001101110000";
            uut_xb <= "111111111100000000110110111";
            uut_yb <= "000000000001011110001101001";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "000000000111000111011010011" OR uut_h_0_1 /= "111111111001011111000001110" OR uut_h_0_2 /= "111111111001111010011101011" OR uut_h_1_0 /= "111111110011000010110011011" OR uut_h_1_1 /= "000000000011001001110110110" OR uut_h_1_2 /= "111111101010100100110010000" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1011100";
              state <= "1100111";
            ELSE
              state <= "1100000";
            END IF;
            uut_rst <= '0';
          WHEN "1100000" =>
            uut_h_0_0_i <= "111111110011100100101101111";
            uut_h_0_1_i <= "000000001100111110010010000";
            uut_h_0_2_i <= "111111111010001000001001011";
            uut_h_1_0_i <= "000000001100111100010101110";
            uut_h_1_1_i <= "000000000100001011010111110";
            uut_h_1_2_i <= "111111110011100101000111000";
            uut_xb <= "111111110001111100010101010";
            uut_yb <= "000000000101100100010101110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110110111000011111100" OR uut_h_0_1 /= "111111111101001111000101111" OR uut_h_0_2 /= "000000001111101101100010110" OR uut_h_1_0 /= "111111111011000100110101010" OR uut_h_1_1 /= "111111110001110010001011100" OR uut_h_1_2 /= "000000010001100011000111100" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1011101";
              state <= "1100111";
            ELSE
              state <= "1100001";
            END IF;
            uut_rst <= '0';
          WHEN "1100001" =>
            uut_h_0_0_i <= "111111111111010001110010111";
            uut_h_0_1_i <= "000000000110100111111111100";
            uut_h_0_2_i <= "111111111001111101100010111";
            uut_h_1_0_i <= "111111111001110001110000011";
            uut_h_1_1_i <= "000000001010000010010001100";
            uut_h_1_2_i <= "111111111011000010100000110";
            uut_xb <= "000000001011100011011110011";
            uut_yb <= "000000001000011000000111111";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110001101111010111111" OR uut_h_0_1 /= "111111111111010110011111101" OR uut_h_0_2 /= "000000010101111010110010110" OR uut_h_1_0 /= "111111111000010100100000100" OR uut_h_1_1 /= "111111110110010110110101100" OR uut_h_1_2 /= "000000000010000001011010110" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1011110";
              state <= "1100111";
            ELSE
              state <= "1100010";
            END IF;
            uut_rst <= '0';
          WHEN "1100010" =>
            uut_h_0_0_i <= "000000001100000001101101110";
            uut_h_0_1_i <= "000000001011001101010000100";
            uut_h_0_2_i <= "000000001100000000000010000";
            uut_h_1_0_i <= "000000001011111000010010100";
            uut_h_1_1_i <= "000000001110101101001111001";
            uut_h_1_2_i <= "111111110010001010000100000";
            uut_xb <= "111111111010010111101111111";
            uut_yb <= "000000000100011111011011100";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111111110110010111101110" OR uut_h_0_1 /= "111111110000011101011101100" OR uut_h_0_2 /= "111111111011011010100100100" OR uut_h_1_0 /= "000000000110101000100000110" OR uut_h_1_1 /= "111111110010011000110111010" OR uut_h_1_2 /= "000000010010000001110101110" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1011111";
              state <= "1100111";
            ELSE
              state <= "1100011";
            END IF;
            uut_rst <= '0';
          WHEN "1100011" =>
            uut_h_0_0_i <= "000000001100001001101110101";
            uut_h_0_1_i <= "111111110101011000001111011";
            uut_h_0_2_i <= "000000000110110110000110000";
            uut_h_1_0_i <= "111111111011111101001101011";
            uut_h_1_1_i <= "000000000000101000011001010";
            uut_h_1_2_i <= "111111111001110011011111111";
            uut_xb <= "000000001101010011111110011";
            uut_yb <= "000000000011101011100101110";
            uut_input_valid <= '1';
            IF uut_h_0_0 /= "111111110011100100101101111" OR uut_h_0_1 /= "000000001100111110010010000" OR uut_h_0_2 /= "111111011100101000110101001" OR uut_h_1_0 /= "000000001100111100010101110" OR uut_h_1_1 /= "000000000100001011010111110" OR uut_h_1_2 /= "000000000011000100001011001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1100000";
              state <= "1100111";
            ELSE
              state <= "1100100";
            END IF;
            uut_rst <= '0';
          WHEN "1100100" =>
            IF uut_h_0_0 /= "111111111111010001110010111" OR uut_h_0_1 /= "000000000110100111111111100" OR uut_h_0_2 /= "000000000010100100011001111" OR uut_h_1_0 /= "111111111001110001110000011" OR uut_h_1_1 /= "000000001010000010010001100" OR uut_h_1_2 /= "000000000010101001111101011" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1100001";
              state <= "1100111";
            ELSE
              state <= "1100101";
            END IF;
            uut_rst <= '0';
          WHEN "1100101" =>
            IF uut_h_0_0 /= "000000001100000001101101110" OR uut_h_0_1 /= "000000001011001101010000100" OR uut_h_0_2 /= "000000000111011101001111101" OR uut_h_1_0 /= "000000001011111000010010100" OR uut_h_1_1 /= "000000001110101101001111001" OR uut_h_1_2 /= "111111110110101100110001011" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1100010";
              state <= "1100111";
            ELSE
              state <= "1100110";
            END IF;
            uut_rst <= '0';
          WHEN "1100110" =>
            IF uut_h_0_0 /= "000000001100001001101110101" OR uut_h_0_1 /= "111111110101011000001111011" OR uut_h_0_2 /= "000000001100011111011000110" OR uut_h_1_0 /= "111111111011111101001101011" OR uut_h_1_1 /= "000000000000101000011001010" OR uut_h_1_2 /= "000000000000101101000111001" OR uut_output_valid /= '1' THEN
              FAIL <= '1';
              FAIL_NUM <= "1100011";
              state <= "1100111";
            ELSE
              state <= "1100111";
            END IF;
            uut_rst <= '0';
          WHEN OTHERS =>
            DONE <= '1';
            uut_rst <= '1';
        END CASE;
      END IF;
    END IF;
  END PROCESS;
END;
