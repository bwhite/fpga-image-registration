/home/brandyn/fpga-image-registration/modules/./smooth_stage/smooth_stage.vhd