/home/brandyn/fpga-image-registration/modules/./vga_input_test/i2c_core.vhd