/home/brandyn/fpga-image-registration/modules/./demo_low_level/demo_low_level_tld.vhd