/home/brandyn/fpga-image-registration/modules/./signed_norm_mult/signed_norm_mult.vhd